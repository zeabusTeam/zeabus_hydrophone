`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SzSecelD6f7LmkryJTwYZaIAS5S0sQmdCutNOKt9Q4f3TfI4nKuaylF8K8IzM3AWFQynyXEhGT1P
KoSsQnB0Ng==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Om7W5npTdDGPn5rJcTLqk2yMupu7TOhcujk5CMD/VPts5d9Si49YmFlV4oTJGGvYm3jZSe9p4VCr
FafDzyEmpR2xbtsu62M6tjVwacoAQWqOHqfrno6N1ZjOKYO432H8auoFcQZQ3xQcy7ZJsiLnYCwP
mCz9/O+odErXMBMcPw4=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mwamp6rhU5u3QyE2cN2AcDE8SqH698UN0LR/AjaVZGEONr/nYNXFglQIVdSfwWUyVN7k+GrSa8NU
v0fo0LnP16qFXLxaCuVnYy4eqHlNoGlE6/Scr5L1MA0wwGVPvSb0YazgXAmhfeam1C44Mlf7uetZ
jpGb5yzUkAPqrmBdnS773Fp2bu5Y3gRPun0ohwRwHPkv1l6/g6qQNvYoL9axqDHs+P3nFjXl6VSx
6zrh1IjAosIouRbs3UbJXbj5CZM9qbuFEkiC645kWPvYWRNxbIg0nvJrtG4agKxl/cp1iwaKHr/i
dZeE56fW5PIhbBrTRWGCQjo4+l5xywPCtdYegg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L7lYzhw+r7nb7cOX28Eytd1anu4DMCUwjrhQaEgcr7/T0n8QUVaan6Fr7WQvFDedIFq4XuBDKhOA
kIo6b05GFlN3ZRc8eCYhbePHFV5c18TofK9NPm02UNIY4WgRxIy7I7TSj53SyeXWBOTow4JJoTDs
S3Q5tU7pUKEUbcs2WNR/pycss3Sny1atkHqahyu6NA/ILs9el+c2P+bvL2Q10nj9WPGELNZSPsmw
E/+XBN8oZccQuaBvbY/q0mAZE/Yw2TzvcurVJL9jZWdVFJxOYkHt1KIOKMxZuLgg+aCHO04SMmtA
70VcXPXe0VKxf7OxDsyL3k6HcooS+k/ylAjM3A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RVrM0WJjwvJPp2A1BBLI9ExIZKJlykA97DJn/U3JtmM5BcuORiNwmDgiJhwiPtKULRkW6QJmKiYs
FTFb0t6FCd9BnaPvC4gvDwFim6gHgoMcmHySSpyyy3rteYOsYnkjcs0tjEKItPV9+yzkPx1a+fAA
m5jYv0V46niHxHh8rSZSXoq2hAvOJeuWDxpr4ko3+tiz1VhWBjFIHLzEz+raaw0nMitUJIED1h7R
kPx2hSHO6jnsia46ABL1Ixuf+AQ7UXZ6f2yoDQdo6AfRmpYgIIc3mmjcRfoYRbgkiFGpwYbQCv+I
5vHKZDjhW16cG1kBH0WtHZOdNLY2Odip4l3qig==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FoQveUWOC83S8UPpluGsTYrLvYhiSMgKuZgP6j2C8ecIT+YpF2vaka4jqh84uUOzaMRZ78SBAB/E
EWDiyAt9l7GjLJm8w89C2Ca9YfHjU00l6kMWrT8Olk5WdgsBZizeT3lY71WQJB6zYo2If5tkJRXV
VzpnE0YejFBjp7L7UTk=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F5wSzisUZZWcIyLjjZYP53S2M4XLAfxlRaBRF//m5y944mV+HeZ6kxDrZCFlneaAHH+gSpF3a9mI
RGmr4hjfhgNrXMwpdLwhKZc/rtUndjoFH6G/GpDVVrJYDpNXA4SSAQp7Bc8V4G4679yxQ2VcyDBG
xUeDpTk+jN1kNI/4MMY/7R4ZBQGuMwBDUz5udteD2m0ut8fFwFkcFVUACdVvIedzNrqcdT4ja7Uj
iCbADUyFHyaNXcoclOuDDNsG6M/tyLpRtU2mwcrg5jBrVo2sb/hE3/jcHuv8Es+pE6FAn8eW6Yrg
4vKjZYhMYVAqkToYafH+DfoDXBWvSU+VbocFJQ==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WmemOUSRIDoY64LsNltKtFBvehZAbjPMFuEy81UdBMy5cJ5tCuOzlztMxMJbfgw5KTyCUUVvTdWE
lo9iXn8XRcHsvG/kwF+mPOHD+f6L5A0jDMWh/FKRhw8dW3aJg3ovYsy3FrStCwgHprOt12Gw4oQe
YjvMBSSHkGNaDkeVyqtq/Y7AfXIGy2r3+HNTJzzIfKiCkb6o9ZAvQZGAdXofKIrKdRRFz39k0h2c
NlCOIVi62HjYniIq/zhvrmGfviIa+oU+FYa57/NYHbDg9zo15VZ+cViPgoUDtjNy9LmvmjN+8wyP
8bENbFnrPMct4TTPIgsH8+drT9Ylur8gODb5MA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 98368)
`protect data_block
j1EOISzrjvSD9BTydNWVgzaJXnPYbQm8gqZKvyskBKBnB6R2jtvyqV30ef/9YQOITNJNIwxQ4c00
/NlpvmR15KENJqXC1x4JBN91Bz4HOazYC3ovfr8notVyjpadXBZvx7AL/pybEY5g1+rF3rd1VJVW
svXi0GNLztMQJDsVIPK0wGyAz7fePkx6S/BCWs0hylF8jf7IAqyZ1rak3WIMefxtBw8YPCTO41v4
P3Gb90sgncCYQ0tylfF38iJEf3/LN/37KQriph79ArjANVvn8e4dSADHqbFeWwsp4aGDqBuHK2rt
mk2D+GTDfeto4zWYXhUFvGC8nTIzkfFh6A+Aa3r46RbBULE1zlY07nLmKOw+6G6BYd+iVA0pmj7P
IRcP8ExoG8wNZWm+L1q3BOsR+XjWDlkJCi3KdrMy0WkbOJ0849+WCfAmTc8sRQS73OJcN9DGpPDu
zlz+9qFjCLnMZOWMY5lfXKLziD2BR0RsoFOWlyiJl7HOeIjtBFWfow1fjbRqe7roKPYZ9wqQa96f
rhAtdW/gu6eWlc1sAKLzEquV9Pq5dSrKLrdDu9AjxYKr9Yd7TdcWwcvuNXY7iG57JSJSGC8zFc9d
PcV6fhVvGzxsUU9kYZOhH9fzT14KFaqpPB/f41Jv7l4F7v3rmZOHN7W0PHlhmjDEjsNLlRotohz4
povhDq1iCu/3J18o87pyT0TFX90WGAkkhJkqDCSv0BlJyr5V9U7YrutDzLad6H/zzdzimdtcNeu2
YR4G/nssfsxeiKVNaGPAMDOzsLaxbBTKN2jIZARkOT1E+NKj0l2oz7QeTCE0xquv6XvlPF8YiCBV
WWUCraoNuBg6uImFVETAA9/qpNSQthlY+NlviSK52dJNmx+wIgkhoRuln0M5v8DDFGal42Ycwu5Z
aeLDGLde+PQwfNUbfZyjh1eR+TZmEZKF0KXartMiN6fR16XyXTUHE5M6Dk6yo6A60ABHziLUrVAX
SA53e8udxXurcac4vIz/eFJgGnPQuwgNntVmDbxAHg/KzxSzcGP6ZfzVB8pWd8QjQ2kxIUu9Le3/
ZMyclntHc+OJ3YFISIYZqjRHCVnb0H1oW1nn0vgqkuIP1NM4uJLLnz3Lj7X6QNtRmAV5lGazH2t/
a31Xtpgppq8dIewnc4fIx2XocKudkjdno6QNh2knqc/wm2LFilNM0rFxI3BykNHyu+JwRAfjpyD3
j5BKcbnqEcPe1PiZFhA3Fr7yNhuNRYyOWe43uCM6ukandNesILuuLlI+0+N4+AWdfQr/PyR9E4gD
e+dKFyVbqcgUbfXwZGejG4hz6PQ29WPofwzLAOoYmimxTz4EQ6BZnjrwu+3F0G8JowaIQJ4CbAMR
ON8ZIhd7KfEkDsaisEjTrc6qRkkcwMRnf2lDaHdnZCUSEjFJp/jO61OynKC1hgsjVyHr1fcfi2bo
3L/aetAL0PK9oCrIkYPRdE2yz186hNBrkZCQCFAEA2/oIjgckKuum9eQOSf0xUGvuRY9ahGGsrXX
CLE+d6ERoKK/hcGj7tjiSFL9A4Vw7vMoAp5H2TK88DLiCzIOLPNvC56uyjV8udf4iJupR79IuqOE
Rf9pGHgcPNszqtNgTjbVF28hZnZq3ICAVcLcilE3gHwRQtsc50CJSGZzWJ2tXRI9iVN0h3DSEfzC
/a8JZz2UGQis1ch3uOhLT3I+4X1PzCPyXTbEhl559z6pcdUcftVn3CBajsLvRhTc3PnYJN5katDY
Pb90MiClFqYtGtJrRJN78jk78BfE/BdnPJOlqJTswYLVC45DsjtOCqAfJbM5z2GzXy1nZxiHxue9
oB9LBWMvpgAPhSAALput8OndBwcTWQMNM4/UN4UV9m3X0LasNleOSitOnQ5LA1baCn1p8qH0tQ3r
85SNxJi8751a1osBBYt7coiJUcNd6VNd3igore3CoNkZsuZRoWdN24UTkXB722NDrbNsKYzCLHme
nJR6m/UCt08TwKVNrmnzgiH1pjv0k8+MH0RXtQX1q8M+uaklAAmY34py3hpvE0RzUQkrkt5hDu47
bpSGaJWJ5Xq/UrF8ja/ntB5oVItmknIPFbv4Uv7zTuYNITCfYnw5NJ6PQ1tJfi9kbB5Zgus88SDV
RD7K4RCp/xZRLd5Su/PIUS2rdYw7J2bib9iexgx4zYjW3ngrJLHvuUf5BQqVmnH1ZoSR4g4hx99d
Kg9zzL8GJwPWiO1Of3p+WGukEUiCL8yDAP9aF4ui+uIEXNirlCxhWDmzX3YfGnX/kkI+KD/T/ptp
DoQoOIAIlU9gfP1DOuJBFV2G8uLeOGtnEn2LpiGiUfzZz5S9ZgMjCVSEQ1bVOzsy20JI9SEepUZs
EicpX6ZphlOUGTsXS+jimjHt3gkWeGIeS03i169Buz8oL91mezXqsqfO9/kAafQScbNCjw3XzU+b
MOiKTD2kmoKELoVGptqhuKHelFwOyvFYBDFuMHPjdYPBFIbXNbiYlIDzkyvinvcrcB1YWffo+mCI
YMufr5g2EOkFo2trHeX2QxcstTrPyIb8cu86CBRV0sPZ2kW8v9/oE2B5Uzc0b7FcpDqJ+yuGQazI
Lw7RpXgK2ucvMOsRrpZJKJ0VP3v4AcdAFcMdzZ/aFFLnMWAjM/OdWTAL/I2o0bUhCSyI4WCottOI
3/08sLVJmhjoGhVqodoX4KT0YwzRtB9ZoJC/1jomCOz60cXCkY38iUS6QIQp2Q2J8TbQzTHEQvs2
LbgOeUkgcOM6jXWgIY2tgSV16PcV4qq1qp/aVoChsFVyajguf96/NtWolfMmeHynGpYTAX9hkiyc
qJDsYgL4VD7FXnuZWcPXO35SYVr1+JFe/CWUphkj46jy+B1mlkUItasNfA2KaH2ImorB2OY9Ew+6
JzUAcGHjgT+fiS2NFwzau/a0GOV9tsPNdsxicy4R69oJo7vQtM6CI5GKXKuSuU9xBMjAPco6lyGy
aT8FDPZjhUOO8qU8iSA2G8HX8/SpzBK0Pw7mO/DeT/OlOuX97oGpP+lZjk6e65+U1gETF0FVPWMJ
dh0bPAkc3hnZfheyVo0TagRJvSjjtK4tnwQgZbGNBnfhaAB1a5P8Aj6BEpSt12Vu+CLQv5z56Bxo
7ifHrv/DJs2OUT2Ex/ttHVbz74iYxPnYHoH0SI6oSTEhThpFiSedsC/vJvdFEEMlCASS0HOnb8EY
+ODp2TjmApb57fvUzZ3t6n/7l8vuthjpfct9Lv7mQmMQ7K7X5bQAydCHd21dqJtUkRSHnxwLZyb0
kVajqWoXdpJepkB1jnFmWCPyRYlTw3/EwbV6OTiNnOAN8ErVdpKKEeAgLZ6/e3zXaH+Yl+e7VdIa
QCpK83Kj8gKdqGKG7FWRdKTcerbjOduiZ2I1X9yJOAIJT7tJjf6GPY2aYA+lVrSw7vZIfFKmCeog
Kxxrp6o4LvvJEyZj9ZW6+HcbTdMcqw7PbbsaCouywYhH7s7VjcuOQ/bPPe/+E8+rlih53K044Yfm
uWy5z358ojfTL4WWG8Mx9qI8+f6s+NwgOH0k4zcetFTd69s4jzolsUmpU6oJhevVPRvHgiXtZdNs
y5mwBUlBrdH2qeo5koKmHBjZfn1Etj6shOsMRuFihIhbY41+s7BiebtnGoql07XwELFDyssseog0
cczy4DMIO8brslveOdR4T0PzI44lqwiDHWIDYBUlpeylrNb/FhXLVv9lkny63/cH6rY3H8+9umJb
c4xv9w9tTTtmVRtqinlmVXQ545NpjdqFNs7ZkZUcZUMf6H8gFFDCSXALBxcp/19XcyBcTvfOhgN2
2dvXmNy58jMDxOqGUg/suhGAwU4gi0gE3mY0C5p7KllAEnL+4kSFgJch5o4/3sE8+AUYKWlXhROx
xeLDfLejGBjVrVfvhAzIk4GUGVeXcPztY/FA+N4mQu0WYXrqScAjBgZ4klTdRrw5+pARZthpaPle
kACJsrTokPkKXgkpc1EGcH3ph0rXkKHp0U9sAYQ2DmZ0Gxbh7FgVS190IfPEEtC3MFe4SClCWZdF
yozQL/oDdj+QPg+aiYwo1Ksn+Z6PMCiYkdwmwYbLPydusuLr4x5ujVRmDZIweKtHgD7hxEmbSwgV
FEASH34hs3gU/Z00sMpP/sJYX1sS3UsB0ycoWdJZTtiaRnuXYJpi7ZFnW7QKRahbkfWRP83E5+5U
QszVxGLSww21Ry2ay0L75xvJOYJ667vGSeax7A2IUMgcNSyrB0kw/n3vBeb3u/7XOFtLs50Z+CN6
CFqaF+7Gw9/0cSI/5pEGy2hm1K/X9dAFP2XSr8Dzdbv7hyVseVyfHXfTK186+xZQglMN6QPjLO5E
8B+J7qd9ro99OmqrNO9SDLzYZkfQYGcMI1n0oix5h/8uODjMebViS4PfHaZIE4KHSPFmJLz9KEoL
sTcFXKNZ0xuEgG09pROY+hlI9ZwBYOavAb1lH9sux1SoRux6iovN0rXao8tKhSVLI0CgMIaqflhi
K6mG3u7FLC9JTfCKRCnTeqFh87m3t2uAaWP6uNe23sgj2bWRXpzzojeUpjl+bmUzQhW1BKRs9Sn8
adpT3jAkDV711ZeWZByBV1aW8C7xbTe1s8yzBidheEopXErSvPS8R6ARRPc0wQfFF3BpACvAnnMM
iDonl3Ltop9L9wOwtZS7Y+Mk3QWKu1ZX+kfEOvInSbyS6FhF88Qi/GFveWdL4siqKwFXbqH9QkUD
JHpPrtZaaH1qRx8/ECOybOY7iPPWOUYEatYwSOBuBglBQOLW5U2LszOQwoxgbHLGU+25zw9OxaKL
6/xqeoZl4bb+nnnC2sCpfehb67W/vBLPfIGWw31Jpw6oCFgenEyoUKHP4CfvgKWiD7q0Oo9OzC5I
0PUKItMna3l4+jlYwEUm5b80L61m2hIUMFvBJt1YqJS3dDuAGDAuZEJN0KE5KSw2gbE6KVxQZ3z+
oSgKaU4XfVA+kCpd9QwZuamiQomDL8KNYT2KlWMA0B97y+WjjpbrOQiMNEHCcZp03MfkonGCgCEK
wd/RF/21vmjpD7Gjad3GQcltCWdM4Gs0jOzpOfNYvl328My9SVnJM0VJ2UUKRypHbYenA18QXDhR
LTkONAV8saCe1ILX202MuukMgaxch/LkteXlEBYZqlpHEmJS9OGYc8h+ztpPGf01tocrgN3RumcT
sk0DP4gSfaKkUP0/XYVy7IfeFGi9I5+uaPaFhvp3y+L+h+80lQp0TA46qf7kHu1GYrV2q4wochG4
dKVOw68UkQ9XrsawReiJrZItBBp3VgQPH31EARf+gV5ubnj0jKZb8QjuLQEtPebo+MsRhTdWe+kG
gPdFRVtbAC7K3IXCqFo2wOsIkbXFTogn0VvXR/Xk6ahSW2q9sG10RVTXzhpr6ItW5hCvMgbFSBd3
YLQXaL5RQ23DaCo1e1ehHmULTWmHvirx59AR9fAEXhhUxA3J4QQW5US6eUyQjVFzxxepexP2JY/9
3Dmz6+CrNbAJd7AbVBDHKeVqQ7ZvibZ12A56SCQx5z3Ny95AlvNhH5WUXi5lwFKOgV08weXmVcjD
KSuGM7vq2+vbVJ8OJxb/DzZI6w2dI7i/iX2HL/yU83KPyP49Zh02ZdXGOkwpGTAWoLLwLUN4Op9N
SDYg35fliGc1e/gN7N/BnhHMIpsor/kYy7saGc8S2kyboQ7xxyV9YHOXoxAp5mg8Qj/MyjLTsfD2
8kHS3VGGi6tkDUN1s0gqaewtKrVlxpk7Bep4ramzIEpM/sr3mTtF3+7CcV2Rst5U04+ZAhvHKJhz
8Uew5lLCQ244zcQ1tskmFFzMU4Rp4bZfpZA+AAmBG1OCfCC9BtbY6oQlkCOtYt9dV+cdcuOIcmVv
fo+W2lKEDq3vOiXTCxCLTiMsDpZBfDLWTCq64ZsbcOvFiaB+y67C5IaELWEYaXfpGm8xHdjiONKS
yO5AfhKBHYHCZKDaxesYZMom+vwOH55RRxLtMYGYiM38qXMRuRnF9rnpmTz8p4mn1vOW/XViw1TL
qpJAFDM0iEahgHqXozyqajpnlljbmAlqvtv7G2HBU83n4l9V8OdMDvEP4M9tg3fCiHnsC+B9+iC9
Sr5MMbQmPVdaAKFs1934NVZHcl3w+lU4K22iecZ2uVEH1Yh2XY8vgO2/anxUWv1poMLa09UUWhLc
9/WqAONANXfqP4HRtflXRUiIL9K6II37lrPr9KuGDh1uuKAZ1+9dFk09fKyE6VfN26wT21VdFvvh
PuAbLPbC1a/30YerFAt7KeuXnB+sQpKS0w+dazbCvfKMt3pCraY+5aRe8TSAIzg+mJ6+d2X5xN6E
BnxOMbi2pYM/0+fOLqfmrydT4qZ6bb3LisH2oH/SlcoQi+zHJ5eW+t9zhggt2KURD0gRXpt+rk88
NUw3tpYJj7c78ddSZciouzAxQxxdMaMv9WZ2ZqhT7yyZlFYXG6sBYd9re2hTKVXBJMRBN97FSFKs
+LPL2qVEa0TTRClhFznG+pbzXC0ZqZNPQ4kfqxyEx9UQGqpzWvYpVS5TIwrX0hLkyJyEkWrMy1xv
gVg59xiayVBZdvOXQb2qxNE+5gzjWuAFtVHqjtqE4lhcytVpqIiAhSgLIwv+QllKibhf6i4z/KGJ
4w8lt6QywpJ8Ny6Myzvr5qiws5g9V0d8Zpvee+//seexC4s0HwGaIDIdgg4aVWVcRMi0m5H5ZzQ4
zk3FbC8fAcsempEhN6iCedpmYL5odGHxz/ldbjeZQUNr4ptBo1nofj4sm55t3Cm79FmIsvBuTY9r
wSRArXLXPoYNGLQm+sSkFZVgXSRy2uldgvUnBurGOTftCXmrvebySHwsxmjjUENH4X95eo6a8ZCt
fsvZ+DnA/lJW3nn2V5fa3/ZZ3xLNhPEZwWuXxK+Rc8SrPoX37H2wmseJkyRKiYo4bDxMYxuTt+0i
rVYysWLZYeNqj3F7QDRBvy5uuB/WrVmqTAi1DnDndnq9eTh+BIAP1jxR2Tnt6at4HgthPcNAfw9E
z6/i/GIcEGA9EY5buIXxhx37ib5urmph/UUjbIuXifcMUvhpFvZOa8wyMb8N2y2RB6VPmKg/ocmz
e9EnkElHj6RWdkmMqtJrMT4Ouq3Zanv+zsJpLi0zszvyHGRbAJMPpCWVBSjlMEkK6RMu2pOrxm/Z
bdtSnvDeBpb6+j0RalJ5SffjjvM0CIWCBv5R/5F9NKLt9G7gHBDpX3nwXTOFIIOzOu06wag3J/0c
dG/szucqIrwEcn574CKnQlLBmeuFfGTvdo5v7SQYkvGfUbbkm1VdG5Tx8oVlVH3DY1uhD6SBNmt7
3AcFEnxLg+kZjHDWCpNBJ67SxJYzKR31dCh9QClYGCU3O/8H8glUnsCG35eLGJbA3VbpdqDv8dKN
hIR4tHFauShpBz7gvyd4Wc/9k/yvmUlEAquJ38rgJvJKQ6QaQoU29izuPLQ46X6cK5OBQUZeA07h
eMZ0jpU/nZXF/l7XCicrdc0a77LPubka/BMuWauk8/GhBSUhCsOmd9YohWo7REDONQgLu35P115L
cBJALkOcAKxS2AH97DLJTostSDTWpkYXlq21Qb/0r+MBbyq6FsNTivSlJmsT1+vPgoUbCwvaf+Wu
zwtlDGdykNmdTBPp+RxikfqTMa05n7b3oktaMYZDb6CkiVHvu5aUfFdQhltgYTQoegIJWnG9i+GI
fsEHScDgILsA++w1dn1GUzvYaNTxcAEN9vNQP5xSn4R7RneR05SUO5zOh6b8mz0IU9pj9u9LFIDi
ZSDuDmcbHVqFtlMswxSmOpFnRAcvFl+wFEgDmP1u9IL+sD2GRVkRJ8I4Tm3sLnWWF3PHWCWNLLeH
IXDTA+I/fMQmxBjieSLZS/5BiyHwW0gSG7lQvS6hpO7KvOtZ0YwHft2zLjoqYSjbIgO78x88eFcB
r3fk1DD+l4iEGpU9DdxeJoeSm6pPoAHUp39IJsbkUVjIxqn+dgLSqAsMOSm8GyYrERXUQuMD34oM
H18Vyw4O/qb6WqVDby2JXx5jY9QDIav2T4fwVeGEjEV2f0SXfP3xU0ajnuTZ5AKL2KnksaqKIwzj
kzFu0QzHKQ334Zt/k7UoUImn0RPAxbBd6ovCsoNK6H15Jsl1ysP/FvduA9a+2ZzMm/UQ1XmPJ3LS
+tcsHuOrHm+JGvVQQbv9ZXB5lnD77ZjnkyZeeH1bLfii4MhUI9FyUCGpTfvbVziDfsTBhmfyX/1S
btqOF9599emaZzufe49f7Q0o9UHnaYGVodzIBLaGM8+ssOOG/IlzGzyYHZnWFsvP9+RMg1CHsPO1
YKEseku1NY/tqihVzeJywPsjB1+hblXp/fiR17MiN3hP4I5XE6bSk9huqtocf/sRf6A1lMcLjoKU
XTFav+NJt8nWzBJf5uyV4JGnbDVdvW1W8dAgGvpAI2mR01XzidTsq4OyDZcWvUayw8dT4vbeliub
yPKa8Ufqg4xdVUiwg6nMH+PGat+O8uGdaGW3+iNCRNueiQZVBlI1DzMBkam88QevWAFgHpWlzoXd
e+jEbQd0KI7vV18CnPFTnfygeu7nvgbc6d7K9wscKmiSHaxP7O8ZIS1hGoUcuwSdfS/6k2W1uQ7M
AsG2zoZpMLxGQlVUTdsNXfwu6FeSpEsG7q5l3FdNMOrTu872GjzfM1pt4qYMRMcQ0t64pFV8etTO
m5cKhWXHm1l6JHqI/D8TCPyrdwBSEkHom2p8Jz+Y12d4b1ukLNoYEHpQNa3ICODJ78WDbv1ABiMp
ddH8kUNSjIrJftgQ9SIoQs/+oe9wePk2HxZQqDd//B0Xq2OdUBFXH52+/pfVwI5PH4xTlFJZ00R9
ti+Hh4uILpScmBOhnxi6xXZy0Pp/ongoyLfBqibuy8eYjIgCr65CQxkUnaMcrwV+ou84sqYDReeq
vJvNpb+dsx2GMjcHAunL2dY6dhqMGs/0epSK69JgqDvw3Hzd4KPcjbMSI23TzS+1YJf63MtblDQ0
ob3kYv559K2jGV1CD90xZfCndE2hKIfGO5U5Q7GiT5VzOm/tRTTWLloZEaTAXDVjV7VEB0alLvu3
VxC4mWBr+GRY+Rvdedt16Uo3FWbN9+HBTlke/8mzr4Iz8RhW5kWoX8R66eWc3C5OdDPt1QVDDuzl
j0WRHOqaMxQluqXrv0OTNuiJvgF+YFv8sZo8ig2d5+wJKfHkfnW/rcOgzXySlkASlae2hgHqAzam
P+YAa/mAMktw0uHMy5kwcqkRb0RvEPDqFTgYHFuxfZXPY41TReDcCP/pSw4MuwSdn2QB7QYiqsle
k+JusTBuPZUlW4NDJw3EQQx+s33FOr5iCfUhLXQ/PF+hdx46zH4hr8Qcyq5F3RgHll6i7/cng8++
qVu+Tb0do9jicfqYzG9L/oxTEgaNVyWuPfFiE1oh+RYCQpWe9FG4U+03Le77CCVD5ay+UImYw8Eg
S3+dihdSyz0U8DetoLagLkPkNwvvToj1Re0UbHYPvivUMDzTjhiSql/OwiakqeYEIjRMzZ+z6mPy
Na/Buzavoo+kjaVGF0ybzjKPgl/Eh2CRd7dcpS2MVkjaPC2HuX0Sy5orI/P/JDUtpWTmbmSkHQtg
A+di1pp6cBshWjwtzJYRidgBiV9bXQ3kXoyVqpio9K4hKYk8nSPIFnJEY5wvdnq6XptWIPX2luL8
PW8PDrJ/4B7scdqSQAiP3QdqWrR9iWPgOPu3zPdoHofWx8J/nYMm+zEdcTuaYndChotPmW5+TKc2
YpJrcsRXkofvDahz5/vknKiMTO4b15ERYZB5wZRMgYBlcp4bGlFYb4my+GfpOmds6h1HsKEHOTwI
aG5jO+L9XhbzVs82bp3DhIzZMOFHaN4tC8oyEUwydl10QGnt+kQf/ztDTsYffCSYL98KlyhVPhJI
wqCP5r0uwveJ6r0ENwx3iZbIGDaDvoN2ci1l9NqQkvF9zORpLXf/DkF8iP4A2joNmXHcVA3pZpMB
jlair0bxMiMV+Xx6oLscsUDPvegxM9+LfQaFidRMfSoz/xTb9sF/KddQKk/8iuBD2eB0dCEzUxs0
65eHpL9F/dMZFIrNRt3AqznQZkT0u5QPjbt9INIEN3f+Chfmifun/5tdH1oXBV2E5U4SOvzMMUwg
cFKDkxT42jYYyi8KyjzJIRgrZcfUqGOSBSnjZoYVqNfj8+ApFfc3H9+/3hd39XMyumZy0vkhejNj
LGEpaETIH0xovJnEa/+Bh6MVtKzmEcYgSxFd4zze68vdFz+N/etGXctIzdlHoGWsKohlISfTHzIf
7M2/AQkXYOdNg64h2ln7a0cbuueoQO6eJa7QyGPKUNwFyFU8B/5nAky0Qdivsqc1cp/50kNzljwS
f4P0cgkqBObl7/3s62TdEIYd8OJzRHxre10AzGbssQxYxIB2C8fEFLMFMyAHbLdWv3tQ64W9GqQ/
Kedw23oHCV79mkigm+cCZigqn4swDdZZ7wzWD9Re+aMhjQu/nrs1lXhqz9ZmAzXEL5SdokWtfGHN
+6tUjBYnFyZ4ybXdmRD/5ZWJVwUqkBd4jPB5VxXngrz+wjBFMpc4UiguJWB0JNxhHDs1ZmDPK/rs
LGm1f6Op4XAfREvU112M+PAjVwBtFLjL+Wie9byEJqz+Z8eSMKxmJ90eXvRFxghj1QzKNmKoNidy
gaYvlveUqiP37roXx3CUbp3oHObsjEBl6Wxu9TbdaCK8MMpcd0NZDr1q1xrfz4BUVyHtepiCKQUq
9xkXh9W0iuRUwSZCFLWV+sQ0YWfJtkg1fikqtcyRGmskNcHbKg65EoygrIFUkcC9zYXlfyedJdqZ
XT6zWjLDed8yoNwPQt7TfQb9pS8BAgI+gDrt6ZGPci/CaC8MME8Ign2ADtej+9nyoANO8TDqv4Po
APfyagEHDqoVV8Q9P4iClbuAtpK9of17xDBpAmsziytzOI5xPNydr9kkku0GpU3Ap3A8Fevvzfiv
J2shCR5W6GklgXoGv0q1kRleH2z/PHQBisk5pDSQHhNRE1wWgYb4z/i+UZ4yQEXLFYhMRNAJa0SG
pxmIFwMQujJZkvUOckpNZNFk9PJf5Z+otrdxXgzexQMUoSpVuxpj2y2Je7O6Kx7iu+pbQw6w+C/K
uW2kcIxcsH4u26WHv7O5otiboH+iOdRcRRVGS1IQ3DuqXISEt3EkwgDdUsbZqsZiuoFbHEz8QNKb
8V2BZdYojCWNIfasOY0YXIMLUFNwmgQJPK/i0fmqedmf7l2kHpmQxMwYKn2F+ERDkfwCS7JfDabU
WNI8swdMcZFAmOWUSm31qLMAeIJd14+BgFr+VsNcyG43Lw51oRf9iaQ/uP76ySxBIcumvgvp2Acf
nUHzzltQgGAndE8M7vSEvaWCVupHrYvlloAFp4EAC2JiW0larF/5XJSVDKxuRAqIx/c7o3kWG8VY
hfc4qz/U721Tz7uS3scXg79u/oDlQCtWADhRHnQS1N3QZFJriW2M7I3wFZtZ61hKFihnJoWGpoua
ZVExfkfd4NZISR5xv+A3o1cAjV7WbQ7ANG2HYoIMjFzj07Eq45fAN4kKhus93qCFRts6+XIBhLpj
jUE7eX22q+SU6Kvd0Hvam4Gf3AABVW3aNmEQwa5uoKhWbwwIHw3a6UCecHGtzZBqt/tKmcwNUKJz
G12gNxUIo/5aCBH59TLPUg/J50tZxAU+4izexAnEEYe1T9eviVJYbh0HnRfLZieaTzcS9K2kosS4
f4f2iq7/uZ6P4w6XnwY2Syw4Mc2Os02h52lAwpBT9hc+Ax+TdTkrnHJg+aB7YkKi5PLZIrODfKZK
3c90A3xYl+kxIXwe892jkVkOPHQlfqKOLvTTcTxr95xqqMRx8z6ikD0kIvHsRHDRTz+rkk9Z5VcO
UBhd6R2okuawo47Z6FQ78cmdCv6uyhAFtjMq6ecuPPcGvEooKPhizeUTudqx61UzdLbdVfODdm+A
Ib4b9SsLixnlZ303m+dRr9+LavOOnL6eU4teqa8mA+eQ/1JmEfS+rPBZjtSUs0StpYit60DryYq7
V+oa/Fdoa4XqGKOPT/VNtPrfOcXMLsF9yOEtOqAnMi3XV51NHbIVXg/y0d+9EMQB5zwJ8jWcihOQ
whpcb0patvemdF2jRP+6+EF7bIJDm95ieQ+JQmvgjN/iiheZInJPmmqbduyXfT2JY4dFhUWMpm3M
RkodG/9wlodmcnTkPxy2wNLvGIe0sj6V1YgINDoDePskrnvICE0Y4vq7En5BcJfkLg1l+Zd7/jkK
VwksO7kcg/j9Ch3jt4p9wlrLPQyjGU9y11CDRXw+/dMtybbEYYK6CBPZEmjxCxvgzPpMFRmsJKpc
Dy/8aSUi07TPJQw4A67ikrVUteFpxAnjA+dehXjCBpLc3jPtwUeZdkuDCPU7DWsk2VHFNuWTQPw2
I8ZqeZdan2wC9j19eareKuSd9OijaC1hKwv266gKCGizMIyhJY2tQ8OMC9FOp2qIYQEL5eiM7Yvs
Am6e6hjQcfFyJKNapQc8qjF25ZtkL50jntep0tefFrudi/hOybyr1lRgdmxMYWriviegssXua2Qj
J888f99+idP9M7xxLflJdJx1I0ICjtLYP6TCZrcEkCLaeuAFy2zw4LyDwJuMCfCNlLDnnFXeLDSq
EJzB/AvOmGJAZRP933on2rOwgy/JgtP6sEbwG69/1++yr/WhnONMUw/6LSQMiS7ub5+CG7FVFV+L
zGRZWW67kS1uP2w0dAJK3mfhFYcnefbVm/bxJIbcFVvUjtrXDCFLAZ+4boqB5OY0wkY8fiFVWSXa
zR30Q/MCXVS0y1dDGvQDOAi6DRtnIq7jCW/2F1yhiZuUL3XuUgl0MM9hQ3U8bTg1Qt1rdg9Y7idt
oDZHom7KI2NYAkyWZjTvOPWjgir/d2VQZs0fJAD1ani33cp71ddG1vYOD50n5LooBmVT9xeCTwwt
we3mIbdqjirM/auP3P/iSkNrZollKmzI1QpouEZsEuSXitMYMW8OyPndwRSqwrOvzXZFSFlaP/+Y
zKsEGkvkQCh7gtuYIr919C7PjNEf/WcFJlrSB1ufNl3COpYdyEQAy7EMMb4zRHJAebOENv/pR83E
pXJVWwntJJyKqu0tMy82zUar90f7BWOTPijq5CTgHX3Kq9Ux0O8EN7Sv4PWY0A3qGYvxjZKJy9cy
UAYWj6fv2sYbu4MQNNwkXv/6hk0KyZ6c5/ox78iCZj8Pj35KVYlYXuNh7T/7lOKgWTfyWLIQq/6m
2EmYfpggtHQm6f5DGTCAU77FgiWWo4AlMoR51B+QQA7SCWWHeXno0Ho86kyS3XNATt5JflHiDyiY
nE1KEg76a6XFNdZNjDGoF76B/dVBbBeC3sqaXHBpR4oRTLa80wEv0ObrIxYpJWJtB22g55Aejobl
X9CiOE0JA57ezBVtYHx6vptQlieQnDRIQY9r1IExO3l5lj1xCewZkRfY3wPxUmzEjN2zI59CQ0/h
cjRs9+3jcB1br+2HgWBv3OElPQkL6b2BdWK+APARFhPZcj+d21mpvlRcKcrgpXMc2DN+K0qnDg79
lmp1jDqx65QV0w26Jh2Mq+IG2UEdLua4BGrdJCa6ogehJCOfwBmfkmZ6TpgVdrKzxhOOc25F6GOo
TZO6iLPxXOKCVV6dHcywTS0GRq0KWgPm2LemHc28RZdhMl0my47RKjHwPUZBOK4p8y3/2FVYeAdi
QkNMatlill3Z0bfZxGo2CH6ue/1OhnIjm1yG9cA/ckHkEDa2+/hxpLDKfGLmDqCXTu7vtwtoPlH6
FV1lUUEChUdEUWerMIxmrYCljQGXZa7+bQkKrvj9wNlJhSs7/GKRrJGkE/TUqax2E/uQUkWM9dmd
+xoK0KzK+D63g70dK6bjvRLFmNIs7PQF+0QDdfnaPcrA/o1/MBlQvvuonpg8szKMnJpdvIzunTVT
mRMEnrmluRPFQEuIZFlwG2IXBIBf9AgKNjYTOuOT9ldufuyL6PVMgi7c7TnXx6yLit6qJEf2Z/ja
MvWeZfDyRJ0MyzhlGbWz43kNhuOvy9qxOfcc1MGs1uUrzgdH8rjMBJwI/e43LqDKvrCnBTLq6tsQ
MujtNvKWE0NenXPjGu/rqnIDQAD/1HSrVE9EWaQ9tKFSZsO9OTU/oVvRLW5nn9dkaS72TkvEtWp3
scB2ElpE8UbJ2NtdHjwRBGnf71TzjHcyDgcCUUTqAM7aUwyIWHQSXncgt5F96NEi7qUb1T2+sgay
gykGi+MeAROghFECbIJS46+c+LcQGE6sRsaXq6HP1nnjzvPrVT1n2PaHyhmsvCRJhcFdHidWnjY5
VxLIVox8Nwsor/v9vwWKmzGT8bw4/Gwoh+aKRbHQHfB/xnX63y06OWSeM3zvvgg5y2DpyFqE8wAz
pk7E3LjwMnIp/yYX1qG6YjXLG6ASZAsf/rjDECABGirZCQd9vCKbn5AVzguoeeISq3tmw9diFMh/
fqoyIEChy0gZtKiJ78aDY5vz7FEWD6fhyBoChz4E+lewebMiz1Z6cUfB8l2RsJaYf3if7aTvcd4E
+SUey6QUA8XjkVR2xJh4bqipV/4HbA8SCTFz1YFDC5qsUs8Vld5KifJE+EsHRPTu7+jcVE69dsNl
4+3WKh/CKoDVLfXoKms60m8mn6xTjdwSy6wF8268bBcPaiIgNMM6uXb3676snERv7UfzSTABjDB/
yL4ppr55bvSYkza93LRsbCVAYqxkk6ldEayXqiB88MObkanFMill/WhidJ6wyNBQ8mSKopggwSGb
mcH9Tlr+ntrSVdOJ0a2KjBMPmyt0sxFqlyzyz6QSMlhiijFtqczIZcTinFk2FQmQI1UbbvBkRc/2
1c9XUq4Pw2LAyIkPu8U7l6pSpPQmGzzT/ESMJMfxUMYqFsli+uLrQO7EQflbKZocFp5zI7q/2OZY
oTr4nN5wlDyUZ5P7Emw43esQ8MwhrpDhh1aEkG/o4Do1JJ+EXlMQF5Yw7WKfIZzqCtJDfO3sDqgu
GZc5b5Gt+/mOXmsFCpcyxbLsBfwOb17fyFI69TY4S6VzWcJRQvJ2r+yu6LLouLWoQUlnxe3q5LZM
C0fRo0bdqry2LUhGNvRW4e8C15WT+pKf/CXt3TQijS1cAQv7oh+cVa42kQsDVcaDAGx042bsARSJ
yGz7+3sgnfIai/SNCnFuuwUtyGJf5kWR252mREwB8iX4QwJH1/rmbqT/SU2J+8C9aTHMFirb+fsi
fQHL9qI0OCwFCuPDtiBZqaTix36UU37SH7oERO7FY+UjyTm9ZdlBz8PTHP7I3U5kNBhnaHwzfekq
n/y+QytC45Uu6jYKtIOXKKkHSFhGYJ/+frDEMcFWe3fIYIcad0jMDTrTHY/BLGD7kmaeQJIsGoJe
QJXgzyRoW23pJhVeCcAFokR5WBLj5v8XZd4Aj1LYmt6F3p2LETh0Wr7j7y4F+/AGyQCDG/1lJE1o
NY8U7p3qEK/ZbwSQtbvByrqzGLUUg5WCAroenkgJXOTllDsIGn99rIurNjrjtAxFGYvAHoCfv7+n
+1vWwGjmQHNgAGUWWbfrigWuNhPIiCSXZ6eaZ1q0FfHmk/bTLlMF8DawHAPu8aoZrjm4HgbnqYH0
W5dKGFXQjXxWj9WFdsNX+OhggXwcLtp11X4ayqzyOmAvlG4oqiCVrKji6zcgdGz/fc6YM0eByGxC
j2RcCoXjaPZbgRgBb1zFb4huKD6BSTw7lQ39ZjETtaX7JjRTTYZNqfCSnFOWGL1+4t+jY/keU7eS
4jWz3BuZJmykxwgFvr558UKsCuoOhUoGOHv/5wTbHo83fcbCgD988tu7hqpPqc6+GTwuH/ltugsd
t1yH1Id5Isya+7xv5W5r0O+41mOejFIOrTXdbY8rJhyXMVdmi76VImcKFL7PIBphm0D4uJaNv1l3
YPx3EiaCcS98BP/Bm4Xtl98iMxRIeDm2cLwVmuKdRu2qj9/BLvgH4Xy/oe0ntu4UhbX0NSP0Ej0b
0GC9+MVUsDo5GY4vDQwCr5IuAn94Diw2HIzBcS1uHSo3C9qITQS0Ug1AqW3WJxi/PS5Waa+epPDr
4bAPq7oaOw1BwlutjQT7KJ3NC7YAXtDMi3V5hA3/5Y4TvGKKscO+U1w/wqszB2JpLsoUKiNFr/7L
PECgm/ixYCw2KJOGFAupDvaZh59YbUEUkpM2ipdJP5jMPV3+/MBFVKSCtMa8m8KqVP2NA0DqtdTU
aeP8MDvYoyhdCkAE8cpkS4l4/37Yt01mGxa/EwnHRwH/C9bIihRRKlxZHyQQNl4Nua93S/q9dWxu
UrLtODA4OozVmw4a1tWT7ybkhJ5GCokyKxbkb4rNsjbSMAGslvpnRLKzVJ7qcrXC5vsupHq45HnN
+dyTHP+QnPjwQcn3SoxbdMAIOXRQ+oWek7HYE0O7Oaa0ME9j2d0Fip0L/LKtaxb+f3yMihZWKLFG
lVG9fLQRzGRUZe+0mNP1/5s8s34sz0F15fvhh88HrfbfsRdwl0481yFw1ZsJp4I2QIdgrcAACUeq
CNeIaypUTRyl6PUEt0LahXnGiN5/BbF0jyiphfM6fPUXyXu3I0d58Er8cCx1oSsjv4OtC4gonAzv
hZVxFIUnLhqsyBH2uKxITPmWiN2Ico1o2tZO8/ZzgHFqHreHYAPOLlN29kBeVCij5GRzPJU391D7
RiY5pbZoDHhYhDgLafNqGjRujdwhSpfdxSXoNE0mFEExaRNtgGl7I6FhhvzAorAZh9flqjQthvTw
EAawNtrjBsQ6tPxuLC13dwUhROQrHk4Fg3j+FtopSIgXHOoSFZNtSOEDPpt7yAHGCEils7EJ7IFo
Z62kXL1BURZr56yqccS/i2wruSG0jsMmD456JBxDHBYmZ2UYEYwLwNd9MOskKHB+VkQzC4A1myD/
4QTq3JhdYygWEenHM5BxSdJ9pQmGONtXzCPUsoTzew2JWecWFnrdg9F7luH+wgxIxQbHIKA34/Kp
D9h0vkMwMOK3Noy5i/b4v9u5wPPqSvkKAfihLeGumOeV7y3Spj4Bw7crHqmKsVuJCpLKL3gtjDOR
ySfBWV6WIqKEFz5J2cbwsJ8yuHmicZ7e+YQBl0GYURnP5ilj1RbGYMEILdiJ49OmjoKRY/RUjy41
dzJKDh8jx3FUFLbjh9UkIfvV8IpNpKccR+KdszcCQBl6OBrzo8oBkG/A6pYpCNba/j1LUavfubSm
13sA/FmoQMARDZWKdnVd3vvj8/Ei69Yic08SGoAfLuHO+eWNtikOHD9TVYX5lPlPi/E2z4DsLLq+
qQmifO5TUziaZyNn9R7ETadaZi16g7drVeUaAuTgf0A6WcR6IbZDEUHutp7xCmEsW4oqOWPEJDU7
CL8Sesdq4fVPO2vjhPu1biMxZhf0uq06WqS1QI4Dc6WBRkpsiCIsYYWIF0AKbR0oVr/i4gip/kMl
4zQTUNUuVT4Dh+/ew8XEzCZrYktDp0rZp5bVHBYpdn+PX336QpHI3erRST3HexUZpgMhRAhiAE69
e+A6Suww9nqGfVUvPSgURIi49upsuoNE7O1JEmxUSRYmhl3kUxjdTHxSDrWkgILE7Z3+wQyg37Hy
bueycRCWUCT+bsn52vqCmEkPHXCKnZhnyClwJiQkDXjQ8gtMOqYb+1UR/HbRsT78w7pzYC86Vtw4
EaLzVcu2h446U78rtkoDnnJRKjcVRf7AB45LJSLl/NlLlGHbfTqnd6Z9Q1h8on7mmDMAzIxCer1C
i2m7qKAuEVcseZvUKUE3EnabxGtVxCcVXReFb8oXqAF0KquSVVIKcD9612s5MpHkWgRckSig9B1Z
/hUGb+X7cWsebx8MhtLmGGYEKSPK+taRROaPDP6oEANXk0/bP9rCwLrI83zP8jckdmVXQoX5RStM
HSAOCe+Wauge9BhMZJ+QbmqD7t/v39di9yiby9nPrPUGYMzWN9gNHVF6wzNL6oX/b9VmSb7fhnXL
sgUoBfQ1SIkgZ2ZOeCstFef7dxl5sfUHE/GtLcG+kEHSeU0s/7f8bZqilXNLvm/9vDhhQtEQSBbw
miMHUfhOpuu3trviBoPZGPN0zq4ir/OEDEi7APoIYilao5ONtYGBx+MhxQpgyP2wMbs9Sr/NNrAr
0EROXrtY0JzmE2qTCbyNSQRPaemBQUL8xokqGmQzqxDbtE/u0nQ3WAcujvTl8otw4VRyKBJDElzY
vE/gxPxqirExBpuh1FpL2bGV1YADUVJVtUj3YWTI8jKj8bkmUevATU0X61fbjbeHrvBNEW2dFCq/
w7CwNXuovgsMHsKnqtIRSqXVGNiA1oSA8zMK5i2ccp4pjq6VhrmZHkn3jabJjTNjdKO36N0eUXb8
saPuaRt29T2eEjTgWRZT913jgH9p8y8NHC7KsUxgolulxGLiFhQRmckd/0scgiDWw7NI278v+vk/
vNLwzp1j8jwgAST/7RBqHtHB31N+F77g2lPKCXUc2gt0umZw/rj6+FFmGajtnE5ufFuzE4QzwdaH
NmVBAmcSuDmZIavVAZ8vttwND2BuWwO9rRDhKWEoVDupwJ3WETZt8Z4gGwB3xcUk6VHN/x6NYJkn
s1XZCj4SowHmIAhWsmGcTbDg27V47gQGXWAJO0a3tiQKd9SYhL04F0ug5Oa44e0GV1e6k6BLWRD+
juwt1SXVj5jN2tFwNAQXGlzAXneuLymRFGXHoIhgWfi6LqkG/Rha2vtE4ATFi/H+vj5MP7K3enr9
o8WQp3475NjeIzlT3mq2x+rZ63dUVnx/wrgCbocMshdlCfKX1na3K3KoInhHxn6E1j2QdEf6xPz2
w3ixyuwQ+AN82mBrBp0lI64/NGDPHZsB25OXs9aY/gYqR7xJKUL8U5znIxmWfR1w5BJJTH9ViWrc
0jYR+ecNL063rEw3iXkT5qYUHV+6t/rAmFxCVg5e5sOoqiRqUk5hBj8xNx6ZDiLqd2zLUce7oiDG
td7fXqlb53RSJrGJGBMR2HqS9Oz11Hud9C0Cqcb6i6SCf9+rvJ72cMEgN8vNYqcHwuD0gGCYeJUE
D9+WjNUq31NXdks61bkFkl1FhTpAjfV0fMX1+OhQ8cmPloWY4mAvHioXCHz0EgxxMzkF/pEoGhdI
a6EZLiPOzSvoyYVcI3vekmxIz8QUsdPSmmhc3G7RuAeEgSb7b53z1Ty1VQ6YALMC1jsxijVod4Eq
052EBoCTf94v7Yy/k4s0D6+forxqB0O+xqNfW/LAMG0w1wjQebH0HpM3Ml+LUDfZlyEQjCkJUBoM
OJ/S687tLWLb/XiCgQQShpfMHia7cRYx0OCbrYdr9meT145h5mlWLTZEsaUd+BI7J0APHF6ERd5o
Nh2c4i9K/EEFnvIYMkxmKnKg8DQGd3BimkkfKeEI3YwNgIMornzZCStDj8ghDBS146CPrQ/kfLqm
0DAcqYK3z+J2uF7kaZY+sJdFRnCHSHew3MCSrdyEUHzJuIzQzqcsfuZ9OFukPvwsAsUwOTM1Tac5
tHWQkrZrsxGcSB8wMW9EPDJmXVsaH5Dx7Vyyb2QrfIOy0gk4DOHeojMWFL50qV6b9FaNyjCs5sFp
6b/SS6BUda1EBSLXXW0y+aT75ASvvtOnQ++yaB/2kxTwpD13ty7ntZAwDzCQA5fK6GmwySxNTQkC
kq+nQDWqG9zFOs7a8PQku/i8ln/4ANeY1NNS0XPRC5wqIv/TzxF0MXwBcBrG4WniUxUIsMN1nQeg
uMRPKPhGkYmcgkoiFvqaC+vl2/BFo+KNXPi8XABMp/5Eofm0mQDQcTGhHp73RheR+seDHePERk5/
9Jqrh9ena76/edaYtgljE0I8iDWjohOoc6a0QgQKWHjaXWdlLCQMNzcvU0xPSYDfIEJ52nvHCrW8
2vQxBdT63SpmCZeJ8mIInToHpP084ezyqLZJhpECt+iG4z3McaPLq9wou0Acd3Ta+15qxiPD+JEx
yOiWM9LIHvz3Org4FMNcGDd8XudcC0O81Zmy2XYdv2OidUJet/NHPIlDhSPBIqIAW4cWLzzFbxUJ
KTroFY6xHVyohxw/mBNYYL8oDT3YDXAbQ/0yTTisw44YwSbZAvSuVAoCRI5yGOZL9A8PB+zbR8D4
lmj4raIC8M1lrcQGWi//IWSO97OZO4JY2GKxuS1ipwUYFD2XGfBk1rKwdJpcHESHKQ+rOxOaq4cW
z/Zhyoc44ZyAceFMA/tIiqfvYrWTALus10QodUddoK/1orOgrnDTMFKj1cF+8aE8MkyWTUQCWhIq
A2EsKOdn/f+YCJ+47CtL746ybvIKhQlCRePTwDVkOJcqeuR7z02do4DnC9oqgqtqjvzc1S9nwQYw
71x87sJTH5q4ft1oyQ6lEp+IHE6uJJb1185vxnqf+FJF1dYFIQ+z3vB6AWKO/q2L1xbPRCDoaJU4
1/J1McnWgJHfmQClg6XkW2vnZ7lV409eKY8XhNsjI3VLt+5ge+uJGVWNjcWO9/XQKZO7rzAENZAh
FB5o/Whv1Sf6lHIVJOOHq8uHX8xcG1u21PzuBj84FtLLCIJetdZIdd4xoavoToegE+rnozLO76sx
NABs2/symkG0A1dzfTBVlFWpOKGKqcvkXHHCFFh+vf3VYNFT7zrDlHuYb21QCLQe/ERhg5veB5DW
obawXCq22llALIgen/SDmE7d1P7gz9zLPBQhdtb5ClpzAxztUuKejpgx0J1yZsqlc2+YjVkqb1fX
BDr5uxFFtNx5uxEMuU8M7W/ySgVga9biWtsi7k/EwIHAIvyeNtuOJB4XN06M787W2SThy7WHjrcd
r5qLvWpNqC0G/hDuHGkpuE+XW6T3ae9fJFKkB1c03NeLGDVhI/W2dMvLGftHftUw2OqFvy7FcurB
dqn0eXqa9atvSMEY544U5QKnGp2KbQSZce/EwfNnoEkkSZqj1kjuoFDt9Y3BpcmK2KaNZuxEoDUK
AAxc6ENmJZAsuyHLw11TPu/0luPAdkvbR9paMJCTVE5CO4+3cZzJYIS33oCUaBK1/El0u0FsgoZj
EeKquOYy0dn01wzYrVBQmHFcUGueg2DLt/zIETyHd7EGzNx+/uEqDmlERFfJrHAXuqUF/MbbdtyH
fPuJLja5E3kEXRbQ7/2XL37hmsG1EUQXIKmLcsJuFjKTgrCspZFrOZMr8Sd5HOLZ3iFa8by+0AzQ
cTePNADSqLR19HjG/hWFFTAPfXAHhgRqE6xy7LZgSoOGBiCzTTlkXCtnfZ9DsTn8SczsLCAtlx94
01Zyv1rp8XG/7gCUk0HNTtOIVi8PB5bHUTnz48FqeML7U8UcjFGne8dFOjMTLAO+zEjk67q+Ingv
a1v0gTF8iNIsPO+yM+DeAd6cjtCT/YVPYn88ifeFmKqT5iFsp+WgyuMGIJLsanlN4g0EAJtetEEX
MFvzNlr30LzhkpDprD7OriEFW3TWkl+u4YKg+s0z+bk2YVYHW2nJd0JfY3tjKKbxOw6xqxJq6nf3
5ypjsZPvsuzTQRyMBckdVZ24YaGNkNn/Y/sZWwVb3fMbEPr6ReG290RGAWjPVh4sbIWYCwSdsL20
IZEaZp0vA1tdMwC85ZA2+J+hHX1bONH+e7nxj7KebPmTd1RH4PsLskfhmiZCgZnlVAMGRqseX/r5
Ez0sno1H/T8W0YXqXqqkEvIXSm2bOwYliDqAcvFaB1u2zh3SRHtICr1vMPJiDj84xgb73YueGSZ0
sitmjQAkPijJa019a5GrSrUMEwuNP8xvuOBQ8DRYcfiyQOoamjOMuzjCG2P2vV/AN/U0UECLlMyC
JrMYLFtJkP0+64Ha9ozKX9rRDHSpOhzVdDQgO+kcZ4Wr3LUKxBSxbWLxMiLdc/dbFsdsybELSs8a
eZxqqFLJtjJd12GM1nt/PorIhaWsUbs1icLbwRj7ZMUMUufK3c13aC2UaqXURzNMJMoZWp0PZ7nH
6/cu7MWwqhgw0X4yQ9iWukjAfdLRA405TnnxgkunRttRNH50N7efnitSq+mB20eQdO+N2zp/3Cl+
9XAH4PP+8QdSJi9RgDWoTRHk14ZorwogLZLBxdOm7NBxAeDMiPkWXFl47XUquXNoSbLm0u9tQHNx
UMHTXXX87dyhsumE0cAcAwCFWqj6B/3dDlOmtst564a8Mz4G9O3c/DqX3mShl7gODI8x01WI0k+i
4vhOPBXYGcqDP+vh9gDyGXHZ8K+rl2xmovcaO7wvpwPmKMdpALgxzgORhg4R7s3IeUWlAt9JXNs8
tOHoOLgrRUsc1Gew1jp2hEnleCC90VKFApXRtApuQArKc9vc4qcqG/M4wo0lLG4v8JTp5xyf0Qi3
SFtHIEDAKJmoiniOMUonMLSlxe61Rb1n2Oa1N12x2THrzO8E5J0MKaroxpY1kvrMX9MuhotJp1S9
V08KVaDuW83HHGhVzN1R8dQTQBBOctEE+QW1x8Xn7aOHUh/9sp+tejLDeH1wXAwYX0YsIHtUqyvV
Y6QEvXyUtAZp5Fg0LDSo4XMajeRa/llGC2ivREYglWeiX5I3AkF9RDCuOI+QuWCaXtt6R23vJEHw
RNQIzKQ4AAwL+lGV8W2nm/NL29idQeS3lO4gKAUGfEUdx+gf/DsuLPIIlZRp3R6C+zj3c3c+92tt
wJjEVS+4nwRFO8OX3TVOX45tNcicV0i7G5noIne/h5HA6jHdXFs/Pt9WCmskd3gZ6YcGv1e95AF6
1tLe7o76e3UQ3lj88BZwWIv2sSJhp4YL16R6hlA0YqBvVLaWhKb7Raas7tVA8yINJ8yM6mdq5rtB
VA0jOiUNEFhqyjKlRBvLX998UJSYncBTny1aGNHV/XFwabImQT0RQ/mECX2KSlY76dR+nqqJbZxr
PCenbgHqzyk+Y+vAdFeyiisxsYR147R+VLGTUr/kMUvEOxDLnr7FrjqQaON+EqRpDcX9D20rrOc2
1Vyzj9Xqg2VGLFuKbuCxMrSnO8fzPx18EAK7dONdjze0BiW6tVrI2qElaim+deYfvUaGw7b5MxD2
/WrCTaRrwCTePbAi64rM/IaJNG85Cie1Vl+ArniOCY7SpsA2iqDz69ov4bu5XDSpYQab9c2p7IhO
zDFoQT9KdoizPC8i40/vYLEt09FolTouIOaPKTQaRIfTs5W2wH+fE0fM9ar5d2cYowK5UVVcuIBe
P+XpCLodvS6Xt4IgNQNejqJcyLLWqsF4cKjzf58PH1afnexiOhIR9QZFtwJmlpGdmOI7TL93qHSI
zT09ielVvqYJxberNrYWWMXbdH0d7GC28HCaxbkDsc51KZzzhmkRYESBZBXa+E6G03B/kiUxlyx1
KS3HL4VrUSxmU+RQ2yg5TYcNSGqBTJ1nbtrDS5oOPQ8XKoyAWEUWPC6jyO5nXtiTRdYInC/f5SV0
NHRVNPsZnt9uHIvAkxmY9dC/XVbOd5VETiK04VrM01dHQ9ApSM2NuGCJnH68iYZOLjRhjvwYi5JO
bCWm/TwvuprvELLytrpacDwjGkiweu3BTIRdD03kNL2JK2LOWCVfaQjmB9XeCVix4Wc/4N2Fxru+
3/+G11oVkM0Xn1l0oAem6gseoD8yYA4DN+79MhStKwN9kd4lt55FykC1cm6sKZy9EKz473EmkQBo
mWMKnyEsHYGLmlRut384w+YXLwlkpYONbyR1Ag2KimWWOJ2UYlUhvsx2szKetJJt6E9qk9WgZQVM
tC2qH+Mb2IPnlv7zgqbud+nKOD+/QJeT7jBYDqDXl2+ZxZhihaHqrKctW1xH0DQkDz0Yq5XjvOWg
PgQ8LQWSNLLb4pirPBKIBp7RIcJQsbkdBXF+3TOvqJiRyl9resjVCbUhAAknTC0dwmVzhxPqOdoP
IpaUSLfpYzpPjvbSxUb/yl6y9pyXkfacFH7Key2MWQPA8y3nwEb4Il/E8K9fDI+DSgr8AjdzyKnc
nn+UoPj42KZe6m45REFosu+RntBn4m3cLMk9c/4k5fiQKRLNODiKQNohRWBOyrie3Q71XyisiDej
LQZb8GUamansqS1Q+x+fjYimWJDfd6UQp348pRwrpOdu20xjuSMTx8yYdFWjMupTPaFECsYLLM/a
+eGaLyUQmjKGh0nQ3ZteTQApRZFtjr51W6wm+spgO1dk+869iVfr6FFlcMREsFNXAPE9uoIXteK9
CYXaXHdeO7yDz5XXcDxc9PzT5OebJzzB32sH6I7mgWWqlJEhtmD9VUqiHpffmTh8Bo6pETTSEmli
omtWUK/R9xaM6J/yqgLGbL4dXmYhzcYTgrRP85EnGZBpNFQCiVJTbj08r8QMMBGlMjR07cqtwLw9
ptRB3A+wcSuaGwCV6pYX6Cp+yFMkizaJzqk/wg5fB45r1Tz6TgP05M9lLEJ+co56ny2kDdMy7GyT
nvBCu7xnZ1lU71gQIuUJ0shMCBLtDEbpxOGhkbKEvXCgNt81DcXxu6hLXeBNOqcVsyQTJUmDxD4r
QN02bZ2u2jX5dS/7vphmNwqphycJTyx0eBbBEMayP1sO1mSCwiSKeN7Sx3KftQ+tTbn4kGO5BGvb
kbuPHUkObdCBi6qa+5O95j4v6kHG9dQaqe/MWClZNYC7cZfbMayYqqSKFPhW5r4WOuwLaNQEqZyN
60T9UgdISs59E61hUIBjIPIWyBxN6dyc1TEsc8hqhJqD5zWPTK8iU7RNWkRVi0g41wZanJq1//qc
R6XiswVess2fKWOVGQ3+A1OJH8fB9bn+umSd2f9jKrFbXOMT2W9dtrOSYIU+8JSVUDi/s/bNg/2t
1lnWMIEIupoLQMkWKHstr05dNxyeGyscaxstJvDpa9HkZjoQJqXcM8iwQ8Rw6l0OU5+2jyY2Ps1I
kT3JLyuuT5A3XFhu8+l8AscMqm4TOcidWYUoPragRlrJmQ/J3bSYo00w96wWMD7VizE758vXLvJZ
fbQMM8xkQ65e/5KlG2pHMPM/2lb6J0fk1YLSwDiTol5XCewcDBfqI38pmPtT24h48BBdrQmY0pFq
52PmaYaIHdoFGkM8pXAVszRUMLJOlYrV0T0bTLBJFay0+Q9l9RLFd832KopNd8ShRGA+hQqLHH93
vdvLmAvIgOW2szn+McZCYV6uHhrNCDn8S+No8h3nkEfatje1/WnrjsCtRHeaMQOaV4Mb7kIDMHsh
SZUyKsFLt+arl2KwExoXobdBwNQ3NO10FCVKhwCtTWb/mBmoMvvm2IQ3bQisrP/0va0/tdKicNgU
CqlFvHgN08nh++1LPlpi/eAignP6L1webCWYrXk42qLsNR6IfbFpzRUYGKe6dyKifn7LHdBjhhiG
fsfGPSBcG8qhBs85X2dsAJoURT0p8H5IdZEdJ0e9sZBjVN6Als5JQB1D5ofedKfI7lbzhxJJe9Rv
k/QojOi6uGxA6nJBgL34/+TuhGvO8JmDHo/VKP7qNMAFbpv7HSZvtnsoArmxEut9mW2Pw/A0a0Kj
BNsDpsTyTLT1RRQ2lwgBO6asbSqjDVSWbRzxkJlF6zVOr27qtNHxoLR8+zjLOpvy5NXldh8wU/j5
nZ4QN2HhAX3nDwsIDmA7hKxV5w9CM89wXFRRjqMq2n2IlbL6URj3h/RuwcHoW/kvSuLZfHE1LTRO
WJjRfAJyW87DuzcayhMoaZ8arFfvbiTia+0lhRmD48wKI1KRgr7pWXQo9nFHnELe3G/Q2E1p5QJ5
oiFBwOMgCCdQYGa3jwDQTBmxU69M07uMLiz7I3qkM3K1OpU30qzbhHns6CkiSPnZI1ie4vIMZmgR
4TwOg6oRJeVYsY8VLYAyeBCJwBB7WWEygmqMjRfA1P+u8mmRO/SPuREAF4N/Tkp9JsxRFSpyYIZN
qTG+9EhYOvmOIKCc6RMWj5Wy61P8FmzIWwm58w48FmRyh5K/ErDiBqlhaky3mjgeBksfLQ9QLeF1
tkNp5cAM46T3C9QUuOiy0MfNMTw+oXjQbuo+tgvjn3eMVWrG4FaY7mCm7kRYzPQSjQcF/JGfNApm
ru0hx/DP5dJjaUjULHm4CX9HH7tSTGa5Yx7oNf7C5WvRe/44vFEP2fLBj+ZzC3ongtmvpX0+9PXT
BTOktHrGNV2ci9NfegwaC9iXX2KZS4YOeFi+ZcnwfH9hGnSKpW6hHaXem8LpzzbiNSWjGnHGzU74
5/6i7QPx3q5u5tlM4n7WqLQRxJlCvxuSGTJMH4dPlP7IUqsazV+rYpRiKS1O0TxwwjFenCB5qEuD
Kenrom5iEX+64zQ3TC5BJM2W6Wq4u3wIinTwtwt6UA3LM9y70lU0PK5oXI6lflwIF2mp/3VxSnPS
uMJqWHMCSV8HB6sXzebgf1P8YQGUSMMH83O2qIY5MeLrF/BOJmm/Xfg2bf1klcuqzwyuheJgS3Dz
fiXxYj76Kn4Crm3x4kfotfy1HfTOHUHXx6V5e+uU0Re5FIaO7BpfXVHa2XSy6J5doPngzkqVrMc+
kez1T3T9agee7L78VpNFhZPAlcX5UpMvR4r6SMSswZMJ7EMc8/0aT744acbbkMVwgv9usB5XqmuD
nllAogEMobHMRpcn+lGI23Dnd6qWfPnHONtLvo4HXSN8tb4tzRwZfCFOMdfX525OvjXfpihP1+Ei
hcck8kLCApSrA9RumJokE7Bt4ogTDbOH0nAb+iWXtsBObF9/urUQFS1dKQA1EMWbRGOp2twG5Ddg
HNXSz3XOqZT5aS/tqKimHucuTGYz9n05pDdDphM05zYMlUCA9PFm1CTusQzw9kALqBVY2us2+tyi
dyjHWd5Xd7c0Lp8OCZ4VX95Vy2iNNeq5Hl55UzxgFw/oI8DZaaRPHiJx+oM5ucj0FqKjXA62eVjR
L6umN2guLQlB8DgNcmf3IrXRWjVzUYyYlGBMEKlN+Jq37aYBEMtXNuj0xq5E/TvuKKujnaaw5HU5
TJqMU2CqUYACvjEFYwCT3IdQxz9ga5yy4GvkLXqLRnCfqrA2GXBmf7ShyDA8C0RSU5PvBIKR369o
UWO6gNRsjWLcq8e3YGDKh+xkQYnBNCCZfmqOR+HCGGDhlCd+JgEeaX5kTnMoY2kXGhwoiiuNzsGi
5AmcWKY6heyArLkIdh9x5u0nVSrWHPr3wT25mL7HQgrxwJUf4EmOeXpaHoLR0Ce53GX7cRR0vhYn
Y17BBTMyuQy9ISaPmb35+1qy5W4sa4ypjC2/e3siO0DESBqpRzwJdDK2QwSJSuiQRrY6WsWrv/R8
GgYJrVS1t8uOeLZ3frJw2muVXuphCNde2ZbbBj1ow7F+qdtsuRT2oWkt7iaHNyEqiXajBTP+DqhU
znfhAYvqLXl4PsMObHmcKJSCSPMsViPkzf3B8lgce7H3gW9S0BG0x2DXITMi2Y1wt8EPF2Oylkkm
8SRA1/w3RC5vDW53UZDxU28sku7Pt6MyWhiO8XRzGj7sprud+DIvPzNUFJTxGDInUJYWxrYxJsAx
zu2+ySk/Jx0jnI4EJPsJqn8SJTGxFLRq3p0M4D8pYBRTg8iNFapiVKXa+IVNjVb7yONko4xkwy1A
n5JTsaAGaj/106eAFBp7v0SxQBk7NfTactg0kvFs/Oek61hQkOGTOtPRPDHazlaOR9+BR2OkRyOf
VqBlThEjwDIF4TQm9R5o0VTB+g5yQhFHibIKIO8jYkOkJuNWreFcaszLYkJTh0+UQUdvbZLBZsxW
wdBIeBM8X6rOivB+rhrib5xcyhoUJpG2zpqgkohFEwZMgtvZdSrWokxN2md2AfPuBqEgnzSdgdh6
XGpVHvf3QcWszY0SJzaEno+P5kdAL2kj6JIJdJe9PLXHNbaCnEM3cefm1jgaxlTRKMMYYkXaIQDf
jtKemS/b0Z/0EGdZ4dOjcCiZEdwzC9ITgi+rlQzwhlMG7jYqcgSYajME7YCsKB/KopQPPbmIdCuq
UJiP7HvY/JMs7owxw3cp99rDPpqL0Sc8iy8WGkwLZEpxwGGzSNkTH5c6Qh0/xT6wouxzA0kL3ksn
DVwGongpu0cQm6+QA092bzagdIxTJwjPcd05XFHlOYhRA7uRFsks7R1QzIl4JRgC03ofNOHPhpom
6+32Sjmj3lVzRie9RW2caf48ckMINt4MruXsWY1ynpMF18qTghy2vCNwOt/2T6ZaPgXkEwbagSz1
Fn9E9fsGnaCv89TadRhHVJUmS4UmFLnA1IamskTdZGwSKzqBWoSh9YAB44FkpEwYvD5/VtrTs4gm
vBa59zsCePQFppXsnvboOQk8cE8UZdQSrDNrrz6SZEJn1iUAEBvOq2Btgcc3kgrobt4Ps4nKM92K
EFg9o202C5quOgSlEAP2uSn0AmqHfNig1F2/v3fPQO1kc9N25N6VHfSQzNQ06MBCk083iqHrcSzg
rh+Td/rBxBD2EhihAJbU8o7lZlAlr/D67KzAU174yxSD1GG7Vo3fsK6I+9RkKu62y9GtVKlXH2LK
D7uUAiNamHIHAxauueigcmXKiwDhm5970I32s4oLswNL7rU5crEgjdJVpfR9ZoULAfatH76Mm/8B
CH7J0WeW8Sw4lQktA1uHn3LjDof9G/+DUONlikQmJml/V44+oWjsqaU6L5+JLk/rHHES54NJiPJy
2zBI8sdCB+KpWPIy8XD6D8sTIxEIttt2WGP/mhYRQ7hK26zT4WbpRaAAZiU3xdV2eZ+1rVrOGhDd
kMycBkluwgfuzkItscEfu6jgXyLJNG8L/tHlMtAmtZ6mNB18BCGWcyrNMrp5DyzDe2TakFVspsdT
XKKKi2JqWdxhjAmJThVIMge6IlhfajlZmsgTONp9KS6Sl3weoeRBZ9btoyonL30vahP9wi2mAu8x
CYXLW20jzef1wdPSGjUYhuODwtt2nTsjdD2VVJyfD/ewyfgbV8Z2jc0eGM+i2kL20GAVZTZALb/x
hFKFwAzuANiTiVspClNS/nVivLT2amyrMlSCKXpGKcqI+UNfx6AAo40zogu1IsQ4sujreSfkhjK1
Gv522oydkC+oT8LZvgZD7IGEP6TLP0Nhw7R2meBJ6GlG3rQgApJpZk5kiPIV8YRXju4DdTEiKCii
R4XuyMb0h2SlENCg+ky++ajDkHMAAM2Rojt/rlqYQnZ73FGY4JRTeev6WZK2SV7v3rP4habRqbVR
rvpCvxSJOlrtemg4tlT6VsEY8C3fTQTTVCz0mwH3SEhyqVpI0+xtatp1Bpo5heZW9b3yPkuzvrEr
I5WKhTKQnDBrJCXKws1wPsSFafTxdIVdObYNZ1Hv/xuuQcJ5MxzfNaA+0advv4iq4rDlVi2Rxr6H
YHWIIkgALYTjRzH7lZRJUmY6RYKpg/X1qh/d5lHYqtaE0LwegACDy9XtXfKOyBXeew4yaf3H5KQl
hsnRalIEmLgpnkSZIDEwhveloUE4lrepPtZwQmNJaZXq4ySI0Djm9za/wdEMLXKsG21Lw1d1NSKb
p7l0FDaijpCT9kp/GGwKnMlnMbQAEyXANH6x0F/btHQXW3jSBBNQiUV2K9j2Lfc1gN7NtH8TuW8N
vEsOPSeX3bmwcXqgA/Etfd5qkWnynKrpXHN/oHvyq9DP7VPAhwU3AJGj3Uwxpy8jvcYdQrEpRtu+
6TyzZUekemKFdVcfBTmOUCOQbv+Hq/P8jVE7z+yP/y3FmRF2LuBwTk2agkpNCI2KPrEVIKOPDhZs
Im0aaEPreJTWfrAAVVqBJL7DIYln/rwWz3x8pAbrhQlvxiWuLc/UbVuQ6CCQnWQrZawyG3k5J5gE
DFAV+2e5RgDr2qe+UQAbCSzNWxP+XBk4cy+/sPjDepU6r8x3i755x+32WkAwKCEZy8E3u832rGvv
TrtrEyOdoKsWGd6ImJ5LAcOX9FWh7i8C14nY/zArEi91i+Trs7/A6rrov5p3xmI8yx62XPf60PqN
6RBGQWqha7RKaVbTdM+w9V0ce0kXqh4HcH3Pn0k/wo0GPn0yzJuJZtKAkL0Yk5Zfyq4uotXhd62b
NBvmhDM2fHXPtFUVZDpAZbnXerZZf0lGMN2GrqCFUrySVwjyjT1O3gNOtwIuOY/3cCZmmnrqf52q
+zCXPXBgdjpbU5y4Now8L/EtL0JH0SgTmDg6/259DestMtEyIWRWsgIl7/XbcN8AFL0CmKvNcj9c
0TSUGB5Y339zufgGDH5i3uu+PwEXU7oIGdc5Su9iBR/+aJy69OKp/vfuouiHieDm7XkUa4wiGibQ
DhLNgIa6Si1TJaIyurScNCd7z59L+0u5S+1hDDA0HWb5poa3+grPAUGOvPpAJTtjxmpKtuxWEkFE
GtJRA6JTrv+mggrMjWAWdVzeJpiFRMVHgBTDzXIEy5AJGgXTDFynYncqWWt4SZQjAz7sIUmJWR1r
oQ4z53B2sGkexdwMWJdTbdN86OUXkK/KoZBbhzZRAAFBicA8ujF8m2bVtgTrB+1hzpNAKPw/j0Lr
sLzIIFd6NbEbTJ9LHXzRBzWQW8w7bxnP0Fw1NDMNnUcfVcRY/0JUyPxHkP9w/B+kEO0NEsf9HgTQ
jNSjwQ4o3Os9Qj/WbS7RSnkTHZHFxOM4VC3e4tDaKaWlXjam6uL/TpiVan0P6u0/QEYxfyF85b83
46c3bLvscQt8z84+6R548x4E6o0c1UaQKAWw5qwRHxsxGwkVpH7554N8+25ssCYGlA4G85XvO1/a
kCI+HhdOd4qpcF1S2f+5B29co58PEREc2wGvVZwagNxaZ0s5cYwiGxuL1ebajl34MZb0i61yId0J
x0LSdkd2zKfi5ROKNQru4nMlXecQ5HX/D2B2hpsVo0rCGYtejRihzwTrlUqGcwS6LHDLPK1mbjxt
LGYNUzvEzQSPm8QEvqlp0PSyDAV9ZdFUxS5NZ6ZksKAqkaejxc8koKxYnSltq7Q/PGNtqQXddWZj
gA1Q+3bKd/UpRWkqquA8B1bXYi71MOnDTh3g58n14t/E+ym0y8nvDDf8jflbzsw/T3kikiC1aoId
5yIcklqJ0kAuXiRCrTMjssZzXK9UTEt86Gv9BUNyb/m8z2ymGp3NydFl93gZfHplpr7xvStMZFgs
I8Ntq1mTs3BA5ygJIF089ZJId5RWmDfyKuDDbTqa3LfPY6mjd3ZOiNUapSWZimthUKXDbMQYYQx5
moOUGMMMaufhvclon/oULlbswRpDhS0Zi7iD43/eZYIAt+oicjRmsJYkAfZLfmctiDylCUbrm8mb
kB9EODJLDD8wnxXge8sWvrHBuv1zbrbOO5Qe6ch0By5t1io9avxt6YuodXPwx1wW80RbyF835Wz2
PW5fAOxdi+ZBRpHhZNr5EhLJPzVr/+CqgYcFJrotYySYWfOs1WBmGXCMgXXpfRfBy3R1dumvN8DU
3ZoYO6xGFj7HmsMX8A+2l1wTWn1IIlLHo/oFKI4PyOqv69UsIn1QaHQvFZ9yR9molzd7yM9VsVfp
zbQqswWL+PAo37E5KZdMp/HQv6HykP20sYE7xi4CF8JoEy9Sag3cw+CQ3H3nkbXkkgfgDbNWxycW
n7Zty2udsS0aibkH+4h24D5R+Bfxu/op2Pe1x/3kHZdhW8M0IXBwxZwYk6v35+caWT3gWiNn0HnJ
rUUDJ0vwFVyeXJn3qtkzHUwrw3yehJw4jNzP4yfrcvDv8yu7uLnZVnO3U8XXn+ogSP/uTor5BFU0
yfIDKVQYlnE93rqk4JMnRd+kQZTxRt71YvLKuX6hLhnu8dyqmXQNayIqUPELCv2tJGplnpgt8YDA
azURQJ+D7POg4xnfShGnyLehIHwg0USGMNHdy6OcShaaQbb5e3G1PctRV0mA18HHob8bdqNa90l5
sPRhtJvy4oSGmeoPrFKVsY6ia+KoSCeTAHh3QrrjdFxk5kzTvgxLArROe03GcS1sGOUTGTEucqhv
FmKNX3OTwXMeTIFQyR75UaU/NhaJmSvoqbviDRQ2c7DtGR90BninzPc7j8UrX1ao6JMYSnULoP9E
2QZwXESn44iTjhoJcTcNCMRgBxTVxEi8eWE9jxMRVhhANo7COqDk7gkkwmMEjsy23LQI/F11LUT6
kqrMplwgA0mQ3f+udSTo7kjiBQb+F3feQ6Mxou9do2H04VA6gLl6a57GRf9gFv6DTwtBVsjGqbOs
LJNg5FwlOMnVRl62S21+BBPHW8gCoaalHN/jlQLhq8LjwsrJu7Kxuq7IoB901vp95Poj1G2G1Icj
BFk9JwRIvCnxhcWmmcyDbsdWhzo0QllONNJpuL2XahQvDXzuZsIFOQSWStmn9n+7LPMJCc6hh8MW
HMaYGckeA6iypnFAcwMC/cfHkk+9lAwjd2YUjNstssKar/pzkWCxC9qgL+n19OWA7O6QqHNu8MiL
V/L3cbdRKcFZ/FoOG8IhkKi3g6cHEVIl1SDikM6+M1Bc7q0oR10XoETHIhWBsT8j1XSQHrp/hwa/
755sr1ObnmctvM2qukV0678PElOnwmPdu8wLLg1vuGtfdvbz+8IVzrWHeWkJJwQ81E5va3YFYnzQ
e3xVEBrc2mG7BKx30qoAYqfgfWCIXAlkNZCiw8KQaXAxQjj2Jw5f3isCxKWOKOmR98YDxlWMokYD
HqIzH12WKXaM3IrVwdNLFBA2pbpcHnQ6i7Cfclur6IMeR8MyCZIUIpcEzJHa1iHb6LMBYsEzOUbt
PpZ9hRD8B0X6RSRFwK11DfcKarufJgW75Ba2jn9qBrlbZyzuLhKSQN7169uRQPwlZWj4XHSOE5A/
4gVt1OTcV18NC7P7q1YjQ9d82ivDK6+A748MY3ok9OsKJIhA3hOIjhQ+O/NsjEqI4ryIH99ne/hm
BNzGZnHgftC65sWy6pPU5GAAjyq+nnlP60LD6PcNcGSMVFfGvByAl8qoJksfz88MPm1doRXQ94HK
EBoYOMgUib0yFWrznAEoPlOOJo3ksiVrfcTemUWBEem34Gdpf7dawimrVYs5esw6gL/mp3l/7lE2
kpX4hEIDfu3hLe0lKP8yvKcH3ZvXC+K0SlLr4LdbdvqQS4CH/btBJ1bFOlMmE1vhFk+qT/PaIT6t
IaunfexHAe1QSu7+Q7M5ZJzJxkWW3U4QOxPsaAUYzlnAp3z3j0vZFF4ho8/prN44Eql2VK4mAwZj
buMBX/tOrNLmYY5XhU47/FJl2gSWlvFFrF9YaZm2pGjfoWzAJPc+EyYJzvQxfsBqAtjLxGVuvtNj
CQJisqbLqM9uZqoQKIlVV9lbUqRNSVfTV578flIHnRbtHABGzHlvz9hDS4BpAvuoqoEJ8iqHtWoV
JamOKzTOAfrMGQAf4K0pw0ltpQmebvcvw7avzOxIj6YrozJCFnMYE3zjRVfwUzp5APlwVZ9/9Ryb
oG66N8QqTWhC9l9ePxZCYsDH2XEcsHGE+neWw0B3v5b6kIfcVzyQPXeG0ia8XT8oez9IUiUgBA2w
kggZHVFoneFHKEZXo15jE7cNSUBPsTcH/uvjnLHegTjgMnb9nwztq5PBFQNZLgmmcJeF9LhEAt+h
CjLmarSy3vTe4CRUEXiyEa7pOn+3EILs0rFxGX4nPP13BJdypDvZhNE2ID9oQDv+sRLPh6LlxY86
Ygk2RZwN8jng0bb7cczay+ydMCfw7VKDApDL7urr1/vVRXrpuFTcDGM0Zd1+K3oDj3UVEmpvhiMt
SOOSRX6PsOiGwHKBnNhKgwmqLDdGXKhwEB4CVYMDjz04EmbmqXfWM6TeM6gcWWAg9+UiA51jGyNs
P0pC+HIBepJLSy1UlcWrUQObUf3ND7t+5QmwiCiXPuFT6CSgJ0EINX0NvfTTHm0VKtiobYtsNeuv
1tMd0O0fCjLcifgZhSi6n9vN25bRgc6uX3oZiCrH+Od3CO643CQWVnz+aZsV6CvC8/zeEC/Qn4bx
yOp+V9geYyVT2JseQw3fZ5ojVmD+Dveckv75vftA8hqQeZn+jLZ+FI/rOGyDeiL/+4lkPo74ikji
sZ6bPvYwjWbrKxaeXT7Wl4rcQytY4U+IpJOjqCx8Jw+7fjHmAiDa7CFvXvUjX9Ba5tpx5Qf724JU
OwwCV8b5OMKJ+QYPGWCatTTsFP1w7ppiV530xphCr/4ZfDQ2rmtVsFimzkX0nh52wD4dGdtSyNDG
6mYlMblwpP0+Ks+11eqDKJuJzhG/vohATMXvmDiv5XBzJEXC0Ulxg+q5cVm8nn6QmJr6BKF9zuyl
u9tEnRCkiDO4QyRKgb07gE3jga+yh3+gMnfiTv9LKvU6CW2dlYIuBitM2Y8DXua4Vv58BpLp8pdw
teADJ0d5y8DviwU3mvisg3+jmLm3roe8A3hzfTtLjPJR7HyTj4rCr6nEfZq24zHwgcH2fgFcXyoZ
ePhYpvfG+Sg1E9mPay9TeQ9B9TBRIdHxFbSfGEzmiBRKqROCs0n9yr/Y8ViSegHn/kYNLe+s0NZR
bOhJDMI+g9XJwnttPOZZIO8TVfr8sVKEC/LawcHmXOqHTUEBlp+VPJQwVOwC7EJrKsz3yWaBQP3t
Tna/pYnxjFLY1Vm+evpk5naF1/bKKjEY6G93HGH4XXWeXsPB4h3u0z5KBWWAfcgKvR4GD3aoOiOA
UB1qzScYhfQ+fqHwi8AJcEi9YvB/NFzKBVMIwXoULAm0SagotTBaN2OFBqyfBVNDtpGTidEpluHz
agknGqqSinPahEtElMv3tO6RlAtP8KBqtDD6o0FQLNh9yAsq38uqbEtkSd02Z4xqLmVE7d8mEEvH
sWlg2kMAdZ7ZzQAqMOlusZJBCQxYlCPu1vrQg531R1tgC6RZ6mtZHfguL+mqkPnhog4exnpVeNCb
w/6ZOY2gqKNL85+O94cVZBphnziMy97GznnbZL4kH3ApDSsNkeRJwJ2XoZZoOBHin3a5tgDGHk5r
MEb5VjWsRhJNtXAJdiaNS/6Nc185dS44XNMfv/rmCw0pwHfWhOzwMOSSnAY+Mh6EGAfADl50U0OS
DHpyeQ6dFhgKpT6RYqpNiO/0kENV1ozuSc4Eg4fYkgz/L3KrHV3L8arnudtN3tcZ3M42ixVmyoFZ
MzkpHJVOT8ReyCdT1D9KA5fAo0Kpx1gvcnXSQqPtp4akEKSM431UPWHcfE3rL7P8faaMyudkqlhe
HULtn6uA71q47f283ipigNBuQ4jF+ofh9e3sD4uI2Wy39bt1ethJmntuU0mHUNdcVbwZg5gdw/04
bg9vleuBb1yOvGBbYAnXDWZHPnQuZ6MUr4nzKszUs3e4cqFV61Eye1r5AvwPIvvRSPsWhKTp0IbU
Bk+wCiVZ6zM4aX4or0nSCYE+f8zgT/CjSxP3Z6eR4gDeAG+OhUpin/wJrYdU4zrfm13l9pD6p96Z
vbsY6lJd42GGf5YTc44AsN3OMiRRTytIHA3cn6V97/VjfYA1Tz6EBLzEAF+yaRFgzIDdFosSQapL
m46CTze5+1dm8wAvEGrNjJobcuxL/UyjmZQGfnYqHDSTxj2X3bUCxcWwksgYjEKFHFQFtD8DbHF7
fgsewjef7R5lZp5cbl6Eteu7r060OBtLM9QW0oWbBjWvm3XMrdk4c9CPK/aw4G5P3sZVsggqxjV+
K2hFK8D65SCuYcoJernAdWXTik2k0lVL6MMo2dgBV0lYCK+6dxmRFFONaQs8DiCehqfTcaxThhTH
ztOk5KZuadSMJPe1ZFr54Ez8t49l2uMw+bZGXXXl4lpPisfWxhc8QEr2vIkEg2Fj+/r2/lPJwS/j
0m1clgU5kaSqOkoemVCSb88/8QduWv8P2ztH0FyzWhjbBwH47dzTChoHlv4IweIDL8Lg0V64zSHZ
ez+VxGc8jcmrsGcqSdXsB6p0EgnKCMJUsgwgKvVjT5XhVkWpgp9Wy+VOVAetoozo2JQOd4mvZDzv
jbBQ8Xkjs2g1ebW6GxsQ4JtL3vlj5dJkQw1LgN+Ax8YkiXf0nS2VNa3Xe0Gi0zuTu9rCM7n3sn74
W9kn5GWWI++gRtSHQp3dQk41fI7+8AwkqkCXRdJA23GzxlBXPuklZT5twtmvCERWqfCOKg23h9BO
NOgVpKp3Vhseejy3rNxMo15rbUfcudtpHUbQXLIGN387rV4RxljwG6X5764wnACTNx7owYivFick
riFZ4z98LKmU9YGauz0kIknH0+M5mtw5kFhCiFN2I5+bnP4Q+7gIX64F1avjZFlVnVbt6A3AVmiC
7AS4mnfeTQzD90kDnMwFjGYpnRlVGpe3UkziL+hsPnlu4QSvYbipyHeA/RVfe/1PX8hcwfeluX0m
RunHaIVb2p8zMjyMqAdED4dyNriPfDRRWzlwJ0hqwYgusDT8I0/LFpt/J85mjksYK1yjDJ9YRMgx
dn8/rwOd5P9zh9MgMwm6ikO2TcMmwNMNOA7hG8Lz2cKFEzsV1VKRPXQcKkr5OrjyaQJ4uEyGgjdG
74XzP5GDCmjQiQYAo1SvZHwiR7LibAhUmK9B59suO9kM0B+y/eQDk1abDbx955Exv/+KlhTpSUuI
zDQDS7pOpMJJdc2Lgcfxe4vwfQnsrLglvVC3xZ/AnutwcJLesxyNzlqPbqpenbk+jVcRQI3vNG6Z
E6L67721o3Mpk+Lkwl7FOkzzcPbtsx8fTiTyNiTRPhky/rlNlfkrL5dvBvfl7jeJon9JTi0v7Rux
rT5MuJx1MR81QCF7JaUKBZgK1n31b4B5dWmrvREM5BDqBU4BjqMxHBUxrMpnkTS36q1OO8+tbyQh
NevuEC72VWdhqkRIs48nm7F9o8R0YVPCSHSbSXyOZzNWPUf9rd8S3zE5sTHrq5iwRZ4XmrtaNjrI
6Gz01Ndz9qf9vlEed4D3mnF+RIWGZNgsJxxpgNT2KV87daNlpGu42H9kZtKQaEPzyV8uvwXUZw2q
R2+I1+W4etOj7bc7yuIf81lp/Hc4wYTUcoB+rGIKVDY3kDb3bjyHh0eOuVyFul/uXXLQbyCMgP/E
iwqHfEForNq7hho5b3FLhJJn5Nus4bJtjvsCGXaXgHHf+dOJF+CfsN4xZwoATDoOinrGxrn6QGXL
C6mQvwNzBxf8s8LPfyZno1YjGkTfLmNiGo0PEUpQkHMg15aaKcq/rxSBxwy0F5xvgo/NcXLdA7zf
Q81jey+8rofJm7t/oIeciK5cX9yIuChAeIRMGdpMFJoeLEy4iLQm8Oj+jo3Knw1UPxEWICOjkxG6
FQzV35BsvKXLHt3ZHjcTzL853INRE5RwbNfsfGt8LABRk+K3Ki5msbdz/YigbCQ6hQWWB22cFYdU
6fzjp6g+q5yp4ioW5fLfo9Lxfk0J2b2c3DvmTzlgTqFBXyLLYvWXeWe8iUWP2sB+7BS3uEzBfBmA
v3yrvs8pzkoPH/ElhTdeY4Y3fUlncSJs9cAAWIpCf3zuywgaTtuqyqeh6koCTIbCEwrpl3FL2hPK
AYdAaCM0Yq8SurxpS3LR+9mR1PXJH8OnV/iYkJzFkyZ1U/7z/viN0wTacIS7XUigCTpFYDM4F4O2
S9iKM9ac9XxA11ioXdAiP6iKUKpPuup/FQCqOW1vuUBDrRAU0BEBxlsgRizXiiES3f3PAliZsAJ5
Rf/H2DDn1NE7A28/TYL+etOrfIUGybf82fAX70tC1nW/w50MrrZCFpxjvQ316N5Un7pHULQmBWQd
J1dtBIy+fzRXeat6AOdE8yu7/8qMJonjCYocGU008Blpqrtiu+qeLNIFQ1agLLuzv9j0wHLiMqrD
5d8zcC+waNBmrvVKLa8jRadexCrvmpyFu0i4225mUMho+4S3YuuXLy3VPek1OCn5Dk/zBTtZPcba
FJR/fxDu/Bn7LP4ygz5PkXKgR41sJ5+VPduUJq36czS61P91jkyufdsyPGs2JPT/2ZfrJbNMxFs8
4ewC8kDPK0PKyYRfqIOQ2FhlP+lA4JpH934SOOcV+YwLsVxj2H1Pa6PVQMHcNmKYs6anu6fj1tXD
tD+iYKT7d1UhPDA3BibR5ZgGY+/D3mJfUMRIfl6ym8TRrrx+sOcwnU5vj+FrIEAJOs2PWBc0esDn
qG7HGfWMijr5x6enimisTcH8bEjBa5sAkL2CXvkaZ1+K9kt2RTzYiaYl4uvKrAcLCrGCrwjDp3Tu
hu8DO53HjfHwJn6wUo7uJ4jwHVsuMAkPqXEQ8aVGUrGmbR/3LhbM7C30L/jMkMNzNbg0KDzSFaXA
TunfHP+H9WTBAyG7LKSiWBRFdn9eGEMzAP2sz3G3Zq7C0F/TJaReaJHx8hsL9sX2N+DXrDCgWEir
K6uvVmBhwYjAxn8wtkUPNjfK2BWdn769hfXkrb+w0w3xtNuo6qp5hIufWBRgLMsNKp4e34Je3Byn
I1XyunRSwvZLibmizXfkKoWWQIUCUwYvOdIiEy6fJEMiKGga4G2nZg0q0QdwuCTVh4wwQ6kA3hi5
kpvA8pmzG7LQ48Bv67vu+ovjdgC/Yus99zzmynmNfj/emAu5bJkYvXWZ0QDypCcOjaw40a+6pUJe
WIfEGXmz/qdPI9RDzQU2yUZ0RmuQ+cYVYLbJReoVbHl/AyndESUvjqcpskQo7a47WoEqpxy2DrVp
16ZwP8l1H1Epv0JZMXXIluDCJyKHac6/bt0w2MCN4lkHPqmSwfJzXjivYKdd5X+bOhnFU0f3mY3N
ZWfrVSmndJJUXacHa6ftXpdKnvI0DATAS90h2iTdI8rllxnqkqArfRyvqvDLBgo4jgIW7pA0CmAI
Ui4kmspYhX6iJUYgnZM+iznfuZjlAfalmun11Q7REfzoJ9iuPFqC8O2sN3JbUfT3YJHx0RI+cdTy
lg2acGUzrH9xzGmdaY2uQaImXsdUrHEiiQVF6R9F0r499qvo4I74PoTVpOudV9qUaq2pEFqA+/2W
sXtHnlr/JXGZa6msa0BABmd8xJ6aGCJ8GxsY2NVcZx3pxq9QOgpOM43XO7BrMtUFHodKqdq8I/Eg
e+EniWPfayW76I9a1yyLA8ifoJyjNo+e7nXsfWpmgcOR9nMCGR42HXIiGkrhpdwtKDOsMOBtWIli
BW8d5aUkv/zEVT/Ceaa/3+37LVVdw3slXZvC3tk1UN2/yBE/V4nxSBy1XKxLks2LLNgp0rB2eBiZ
+K5ZF0AOScV4RBX6atY2F5OAxUggHftEOpwef2ztk7mSEW0Jod1r9v975qx3wFN4s9lNzitRryMf
1jnaxS27HaCXgwtxK1yH0zQ6rm3KQYjKUWGNkGRN/rz/heePUIL6cPznUhzMfZyYldOqvx1qpUnt
qDexTB8zv/UJvT5RWP4+qI2BOoAG6SmxoPsorFCJ0gLFF3LH76k4vEsFxKi0m9lQKxx18KUE54zc
7HP7rw1OlGNmvBAB52C4FI+rT32nex/lPZFS8RIlkH/uvpY5ssYtQ/ZEgoALqrEHS+3JapqduTJL
qeAjgiOqwT/KYOulHXPg1FunvTF0yrqIKUDYtM1thXverXRub92Mzd8HK82ZRlwQbP6k2QeOjBkj
ZYK8dUQIXmHpt9OWopMM/6aNdexuDVU9Wjs7wfUGQUw81rSdDZt6pv65DVpNQZAwK0v/eM5FQNqY
VOpxMOHwI3pGNtxpKJCBgOE9hgTko1z6GvRr5Rg8FI1P6jlelQ/vkNm9eTEnN89deUv1ih/9+VWX
liw2hyaDG+yH0hrR+1wIN1rDYiJZIWbFHcki+UZimswfPDV4oPNHGuhJnj4Uql6PzXcqCmTtFhAs
4A+j9323udnJrlkZZXRv0B8wZLXx3wEwvEkQgf/mP5hOIM2w7glU0nWjdI0vf//JP8S2VRxygtAB
MmU82tuoNLbJ+Jcmyr5xjwSsgPKYE/2gst+v1r/hrYkrGaxeATTKDmcW/PQB9fSYflI8ptuwRsFX
9iLSZrjPYeVCOYOHnaS8+ldYPdUWdxdQucOCE0ctSdnV6YHq0ChCh1HEDzRC7vbHsvkmbMY/cMQV
ruzc93eWV0IQfkq/l/roJlqRJXzE+7ZbAyOIba1LzCooiiNmrGhb+xAZY5LvqUEsEb/ahWV7mZM5
bczIIs+PvWbAasn7RkJayCJ6Gf2YuUwobQsS8gh19cuyXSzQHSmMi3wmvjmsMmOa+WCiY36BNARa
nhceuK1m99BHpDe2WqzTBOnb8elGVrR1CoKBWGuDPslk1beTa7CmXveLxwsQZb2j9JdPprX5/rk3
BipEuxCpm5D4Y1EYP1A94/T1FBVlB4IlmCmJo4zu1EdKG1ERLLPKl32+UeH8Xb6BsIykve+j6Rrg
F7ixXWH8G/nE7ygFzunodJkoIbFj+DWRl00bmCRRM/cEY5PtEY5HKTPMCave11xLzX4CEpk2LBlw
k+GcBX6+0fYIheuTIJuRBklRWabSt8BqU9t3zF3XM1CnTr5+uhFYOSauO8eowjYx0y5kO76FZ+sG
uaLa7k6rk1vm9vdG2BaxAM4g/4HMVjic8AE8w9tueftXajp+hYmvZQRxlKJzf4IuF4ksaBM7RCJn
qtKWjIosIdyqxXsrTTeTnx6GvXUQEIRo08JMZ0hKWtKISw1knnB866NSGeRqelJ92RCt61pvpUyD
pHsmxrmI7gJscnbJSyivodPGKQKcFJnKxqZiFXAEO14oNrMzK/Fwvk3mela1Dt2DvJv83CakVuzj
Hitb6f/JGV3iwp5FCONlUnTeyDadsMhu8kQUYyAk/NCtq1QbYZyVTcT2Hp8xIBeji+IMSq5WDtN5
Aa7KOu7w074ahrIZDnI71mIPiqv6CGkPLsn1myQH2+us5gKnw2O6j7m7MI6cVa3a/L8LeTa8GKD5
9cIQIQQCwqM10oderKaF3DNhGkZ14uXRO59nkNOnK14/2JDcye+4HlMjllP66hnSmqCYSyxBIFbL
N/RS5IO3WIOZkCEWO2+CQ9kwyTbz65g6sReQBkN1DyAd7S5l/dffVHUzhlBD3+IGPNnYnnJaXV3Y
xBW6UhuDZCb/kLRjBvnMhNfqShAZUSMniTYbgAEzauNLUJzvRyEFMZyku+crCVRxKzk9TyVfmi5o
Y1O0QavNFpA+G1PD0va6xmrP/eIyepK4YA3LBXYXcDyViS1JehmVz3g5qbk2SDFu8+iLyZAz93rE
Oh6Pu92SxE1WW90u4VZjcK9iHiqNnUY4g8qOLdQkvhX2D/WuuXh62+maWAZK3u2h6nPdbTAystEN
s0P2J0RtrgkmT0o0oGVTz8C5QISrGon+LZ+XaQ1Vs8f0c3zz7tk1FbiQJpQ12ZS2otbWKVgw0Jpc
Tly60MVmSOq4vcIfOSb1xnM4Yb8kP42kjBA3yOMSWOkwCObedyIMYVzLoPaoeXihkvBFfZ52q2Bc
XulGgr+ujWnMCGGme77454/ogVUmZWEydSybaGGlQ+iKjBUzCgbHk3Xopk9PXnYYK2sbSmnscU1s
NFBIZSznk7m0RikWi/cha225LSZCL6jeKJU2a7gHNDW7okgqn8CgDmqkAYab6SgHeHcFLI3rutHR
4PkNGh3TLZJvmXU7Nw2pTzPqTtwmoy/mnO+qCRuKijfvV1lpgW5eGlc/TI6bvoNl2U5uTJel3vXy
ExD1ZDPH+czO3BTfWQRKM8PN/pAekbEMsZPr9uLbs8yTmdLZwzZEzAE2V0CXpR8PxWLYnBPA9GxB
bqVDxuXzHai7XnmmvQcPcSnr3K1lCaPHS7s3R7NBVlakMSHNu2HHrgzGXFCDbB9Rij9HY/fEj97/
jf4vhWL0T33gTnwDfwpf8DjVu/WvCyZVmtwP0n5nja2fNpZY1soOOLBfiuQXo8+hlHX9OxIKRY10
QevUwWpuGx8+99r8lj87ZQGIQOs/rJWeQ6MSBvMyP1XPuzXSf7ZbMngYuQ3MTFLeOYN7fK2/wyIi
3qlEaUVml+2PHSOfqdckXeNbdyoCxRrRvFsYMhvAjew7BYqfVtgtA6IP5HgDgCNuLvCareDoT0/9
9gYKfuXmyOQo9l4ZLaqI1DVkO7exCpN0cavKVNNZU4Tl5wcbqFJ8rb2HVuMaHjzVU9OQZUP/fPjr
BVPZtqEvkTivAZrYHcom+gSjSytZsSX0gG+2nSHKBmIO1sIG2kOxLgI+GrIuN3Ktapd/iLjPGkRV
sbplYnAluCy9L9T6wK0ClC5vtipZRTVmND8d/mI3IlBNL/PZQBppyVP3owtjDWGFVYQMppbuRb8m
iKeNF10gR2QItRbzdCLr4kS/WBL+pzcGeWILQ0UdS9oB9tdG7MaQV6q2cQwP0RTMrVeJOS7CtoWp
JBI4it7q7SzQUL/G807dAcNmC2O1NFHrRQEAvpu3VA2aZ4akQEaFmNAaiGxqr5vnfI80E7+k2ck1
+biBzG3z/MeM/JKjhybhYok8PHIo0OPwKYjAy0ESMljXrmQEdZx5zUGb/FdoopGz8mZ1CZKQ6LqJ
QjGjy1qGnlFwILf1FQCaPAcL8j8jkbgldPuuAEXfgPUfFyyBorM8gKT0X1Sgx/RMch992mzn6D5E
CdwdoTEw6TbotNbRfywMFzI5vEKeUkfDSQGynn/Bv+rKCwE/8WOyH4U4CvDm3GkQwkYXGb81Qn4X
RqdzWn2tSJdBkDzvH5zAKmmaG/U5DjYtedMIOx3oUkAegtH8WCAzE59VD+mlDE1CqvAHIACd3/jW
eJLpzJm07c2vbulXqLiujsVgIi6f3udPi9YwstSwzJy60c1FIo6Ku2MfSPN/3dIGxVRFxmeFEbhM
L1aUCxckno90PSVKLJJV3DAaSM3JPu8QMB0+ks1YTLmRE0+ieRWWaiNgzUsBUku3qfDAcMr8sd3C
2vkjA39jJV4af5QFhUN7ieBBB1qyv3xZVZcSeJYCB7iCJj+JSGVfLAXEFh8bhjsMgQx4oGudqNjk
Eep9XiXrJtFKLnEX9BFSb3cJtjfxv+SJIIo5v6Al2aLSzzKwA4mNERCZBcpTtsI3j9ZfdY9lQvfC
H3/0Lk9yh5wy9jj9MqQnu0y5U5p3aXEkSGCiWpSEtTY7P25I13A/hQIpdHjxQ3Nw5WwGv6OUBm8P
6s7dzDSTn4gmcrPTxm5NMJyQUkorGa7RI6ZYeXIkKF1OIoEZtZae2SAS8JFrq24CQWrGsopc7UQ/
mGI8hG/UAgl96Vjd/UB9AbXLt61E85kOPXJ1hBx4pWmb3pcxSx2JZMBW0LRYswxTug3z3qe8YaT4
lJJI3uyQqHW+pESOA8TffH67e74S7co/pakJxzsLvnXYGaqyy7+ZzF0Ehx9cAsu222zKbXlFECsm
70r9Kuxq48vfMfGJatF0cS3f4kNWpVjVDCEp/2vPsxrH2pQsmZl9L+9+zYhwF497vBTuOLysIzT2
vnpWi8WkkkK9/Ml+UXovsC2ohjKA+6e5Hs/0QqAfEJF206PPF7pfjrAy+3ejaclfttXaCX+GhCRB
zBPu1szyPlMUporYjzCi54EBPFMQ28WBlDmTPubFB5naIZ+GwWnUkoh4QH/lDZxQPt/+Fq6HNb1H
+v0ErcSZabCneYpKim+NwZFQNzxWcBX8SRLyjG8eUQCJlqBgsrFZEpjz6szSXl8BF4m3NXcNJkxv
ExIZ08eWYevDKjyDuqqI82/Em0dNDntczUCgQJHYYA8kVPhFg1Jv0E0IWsLF8dEr3lCphn6/Js4K
caUTSozJ6mlNfuSVBaY6VFILWOdAE6FSkQv6qLV6UJHfbglRy6xxyaZUiVjkZxYmDh+j0C3UuXES
TAF/dHUxzjD0mTAT//oC62Iiy+bstl1fk8nzB65mcf4eL7PYjAyZ6VdRanafv/buxzOhUZdbxPd2
GTTjoCjKEGECD/kFJglyd/7jh6wdd9RuvDFsSf2OeSZXbXFWhnJFmIYF1wMO9szcTYtAJDfka3Ky
YJdmgQm7NJgnKxrR2r7msr839YpocXDWDJETHFQBS1E7ZVxFkNAqdvN0hHUaC58OieLb/PjDWlaE
qqffaGxPrlh1+hPHp/DUeAjLtoLqt7eyxoxOav0bb6ZxbTKus7QkR21PRM7S7iZvognM7qTxIz0R
vVHFtI8kAVc22oRBrpWuS+Zn+nQt29Mic2+rst0cs4fhhFWy796uMbxMMKFmECOcDhzu1IDtWXi7
loahTFq96ClA03D7/9pFiOOXqGStcyGp3wqdclxVbdlJtxLsn41c+N5Re1v/Ap0sjZpNGUIrHK3H
yVbIgaXsnyLESEOVpuGkGzqSWZQ/NZxq/MYIIYTHgvYfUYJgVy34l+hapLowFAYKS4WbU7UdZhAA
bdTYE8yim/KOGIWPlLw7vJpOoeWKoVvIzBVCHfh/H/paanZfuVwebp2JzAEDekmrOoVImwHjehAx
Dvkb3N1C8dCZrRwToEKFA3VXpJaNYfdWSppyTxslIJuuREM20dxpCQrxLyQfcsKh9sCrvhaMtdpQ
PP8wBGZ4RlPBJtyYyBGZBN7YYMFyJfXy4RXwsdlcPFfYRdKTWQjfmFp5NiwsJ9vj3XIJy1SR+Cza
7BTf4Ea+EkeV7f3zAjybG9PwQuAijgJwZ2dJiwzgow5Y7bI7jCDPCWsCBHGIEtrcgyEFfHcmpxB3
K03GXYdQMUPfvkRUAuEMhUoUqpn9s1eMFSBSXrTewTEVjRjnhYxDDztBiMWosB/wZsEextYX4iG9
MWEvxEUMGTnrGMg7Nd9BJgE0MKC6xs+P99C5OLy/e8Bovq8RSF/7n5XRw2oBnnNkCWTumLje8O1a
E7VDaNIyzhRt+5Ol4dJzApd3zJ3Zrs6F1W5cC1rZSyx1cxD3bTvnT2rkMSxOrFmkjioYU/UaUq2S
d9Fs+EI2x+SgaJHvdgk1J9xG8lTMrl3ggRMtYh/wEFbgivZDxeXvpp9asqMkSp/ix8NROYO7dC5g
k3NsTAQPLrBG+Ne7x4xzESliS72AjGwLJ5XOW/x9fglJE5o9RDu0DoLC+lHQWO1vWbYrWwk+UU5G
c+3uRJKFjNptv5gjwMe/PG1TmWDo4uGyhYfMco/G0yYZYb6kWuQfjlChdXDmMxmg7L8d8Nc2E4Pv
ZPP8WyCx9S9tofixy7iEbPrYUuaM9iObbeXLoe61+nVHTERpLvBkYPm6wWldrmUPLz/zKdWxiome
JSkJNDnAwF+h2S9txbe+jyKGfudP037LQvrcYsglWTsX0bYb2kKn2ZAzbAStfOqANcJV7qB99knO
cjNgbjPs7CVw6KxdvswyTiph/37e9Y0rKVFeBIKSgNsMiH/rmBbY+NzsTwSNMja/oKcvfgk7M9tB
JNii0EbKtjXUDKEjBLpKu9m6t72wyoFUCHRLhxcdY6ev6rC94BbjJ/Rdos0twCjOObSlMeYyLbpV
Ur8HVk5p96foEzLCTGYhjvJVOykrENi+Ghw3tvdWy609M4hsX3lH4818lNPa6Ls8RD+kK/0ersRp
G3Z8498WfaFj6EJdW6iCiCUe2aGVRfCTYKXWVSx8/D7zKSRUozbKVQUIpBjrEEx7mxhWNWt4CBpv
xYIXlTPp26KZqHORWh1Oh4NpOIe+upz+414XznvpboCH6U/ZE278S+MKmd6QwJe++v38DqsYsYXt
JwueAxgzeZ8AwiBa3H933rptuFlBYi//BShoNO3SEB+5y4fudeIzWPuRW8aQZWG/Y0txAiSdCiXh
V3DIV3rBF9rjBEFoM2lTHD9KfHDDJw9N3C24Dqy0lQKJgMqQW1lQj6HVZYcG56h2AHtlcfCKhe8y
J6W0+KkCSG/XN3S6sbFpmjWRSPt/IrsQ5Naj/fFv4LOqzXjNApMjVgCrldw6MOcgqpKSRj13FTnZ
pkxm5hRDUuuEAue6x6Xqk/y3grJg6fO3Q4LGu+ig6SIpN+47biZP1wTMppURZvg36/rq7kzI3Lwa
DZFL+eTg6U0DP8FtFOqVn8/qNIuqfSVlCOMpVxsR61rk7hKYxDmv+AXLXWsC8nbdXNEPHoOuwG7h
xmFpFqeMOvN6fyEJIQwSf7RGJnkI9xKELtK/8cq3DurYzXk1uySXl8ZC+V0mjcoHUGo+eaJElXxo
V8xHeRCTS1Nx87vYSiMD8xNRvIBiQrf1valFiUdk0qh+NhGQgot5aREdy1IICJk/s5g20GGR47/o
+R/UpRZzbEg+tY3yCUR3nLrv6+sidqXvSSHxJkna0FvhQMvMVjaa15kbAW6l1RukAksun2abQPGT
mKWky8chKpk9LU7irNYE0yzseqnnmXe36Cz9TwUuzBbfkAyo+td2NNNUjNMbeDUwtvp/JUneDB0q
J0M+qByh6nQ25w/AVDuapNmeygdmNI6N9rR1PrYw0+Gmdh8szV5YeDRKNZxg3lMFpvuzv5aulBT5
E4qIGZw75YyWbaGy58Zu6Ef2n2VeuCIYtuzUgHMsw8MM1D//GhqdJW8Ce8oWXHigG8beECkkCLxm
onBcKs5Lpj/mW/hkkDIFVi03wQDwovIFCAFcJBJ5Bbwv1xaSpxhdOTVkg5BoLdOtQ5H5n8ynF22R
Cv/j3XD+8VHaDXhqBtQ5Dyavm378rt4f8XfY5jJIRy81U2C0UJSVS7tHc4niN0c2auQQuerIFzFS
nyu89MUHXBUI7jvxMjx3wTjM7gyNySem0tw0K705T0byasYFoGjFukzSnwmqvf5PxxeM5ZISjw0J
gJUk9kPAvH4Djoh14pcpqdMT3efOw7agfzrVxWTf88DVfjPE3lR2OWfX2s1Fd4j239YqBy8M03N4
yIfB6MTOmUQQSL9Cnp2fvWI2HfZT0C3XO6FFRIoSGckdBLhDXsAJeXxFmi+fXpWh437DuOUtMkFq
AhKMvdw6aYuwwWklG19wnYFbTqUeJ3ack29QXDf9nNZhyufOprh+ECZfMHPbOMjjBm8IXWW2c9on
j1VGrk9yDkFqGf+W8ss6/+ALsvg34SuygmW+/0okNpXM1yvqlFDY18m1lLZ+80zUoh9oBWrY0Uwt
sxzZeLGUUTLuVThrNPhSkJGCM2EBuH5OSUXapGkEfm3OShZuMa1b7wD9RMTxECzR2f0rhJOaj+km
JWXRf2W0BPXY05u6twjrgJ5q3Uj9NttsQykQlvRYpK9mVzMhCF4Po/IofO9RuDLfN9twC9VmDMMv
2jwj/lYbgsmtkFzLEhNhi/SQowA1ol9jGOjUYSDPR8Xb7kp9IQEnOsRtARjFV+M8N9yocxlmIZ2J
opRZCDcrX+MHLRbiNNZ16GZCcW5Wj6YLmUUpwyiv6iw8fjrwqL+wvUOfhi8KSaJHQBehLQ56ikzW
WoCcHmSGXeyjCVYwJOCv6kfawlTIEUZQUrn3oenOfp6UArx/6i9Ef0rxzPLQ6IILN1UY2G6f3rDw
gjWT0/Ke5dvy//8s1kMk+jOMGjOZvJ29+uozuh+izGrixOsFWPSCXOJmCHa21XvuIqK3l9T36hss
oQGb/kaBOu6qlFRDrd0JqB4154MBfmh9KB1JhvQJDxoOG9p9iavWRe070TuPs7bfD4Kjp7Tvb+s1
b6FqbHz7xYGyrSaQTH8LDZdCYlK1+nxzxyn58PsK5DfLtrW/9ILql5AIWe3MOGmPW8qa9OKa/ahs
EZ4KgsU5fqgkk3a0p0YD4HTVHrsEADjn1QBAyuStReg9S+DMPNV8zELO6r5pehiH+KI0v/PN82iY
TSGdD4tTkHMVgoKdeeWyDSDNF7fsSduF25nW7IGaPqA8HU4oFQXjTd0pfkrUzvlP7Njzg3r2q3QI
/eSJxQugr6G9VToWSIjpk2ocujmWaTG208Sto1ej6WluM9Kc8CnHxXsoF7alpqFDgqU2KtwiYLJM
JwrZs1x8eWv7T4fIUYdCHSQvQcXtgXoAq3+SbLNp3V9rLmVgAEf9pNatgDxRzTFN7PS+qtgcccTH
wB6m8x+VDyVETkLN83bQYsAD63vFSUvYAi88Y5/YO0UsYcgqmKvY7QcSW/fJvQiIf3cQDLQYM5GV
fRgKfrUR5+P+LMadza+DQIB5wgOVZjiWd7VdFSU82oaQfuQHvkYXS4zFNBf/H3TqxjrpTj3Wt8Vq
FXRdB4xapEdk7HvIWDMHFO7WGNl8IuCWpafjtY+cUrV3z0iBXGs4+MOUjFnceJCWKV6Od7+28uat
w0qJyT9iJaaDUGxm/pdfSX8XwATBJu5fegKaQmd5xxgyPZMm/zRg2HcdpIdPFRDStQCKceETiwPs
/ACIvpNx/IwfAYUVmlzxcU0F0OIA0VaJns6dS1aLg1CXKt4CdTD/j9WZMR82YXEn9u/f9lrCiIdU
s001SdEPVLYaSvB1pL8eCArMFIxDObD103iopPyKbamNbl39ewH/N9c2+gcZiAcrmrHWbKCzlvJi
1wbphbOLFW80JFjZsWovEDeVAR6AHha0P9rfNBzSo2stmoeonF3Jp4222NubWqgzYZHX5j759R0Z
DziCbObxNn+Vlxu4XepAhHWHn3gjWBs/YKhAtuEZNhqd2bw43Z5OQSPWa9KtoRIWHOz8maiFyJSu
c6bBrBi4PWzXdmAIBgNoJA4u2ncpbdAMaAK9z3K92hp6EOkSI9covFo9e4VOElhBQ4NG2Ttb5BXu
zgrJRLUdpf4r6+2BnNUiLHkqWrcTOU/4oNdfQz4P1j1ykY12EC4oBhW3BFtVWCgMxlOgz1/Jz3pK
wXDpt87C3IYnpqVtvoDI+6XgtjjfGgTFIFjJXmB5i8C3ywAq1p7gqYJB0GhFM4ZxmbyfKEHp5Szf
CnQs61juBk5xOsbZAjXs4HJbRPeh6oWqb86ad+kEYt1q/Wd8bV8Qbmhd0fKRhhy43K6WWnRwEawm
QCS65vCcL8TvhRyvr+B3AAmYlSj1UUKCDUcKVV6D5wsaiB29HNj+nBzZ86QmnWs90cmJ2XO4XCky
RwlpHZk5/REQ9rXuG7mYtClJE+MXimZ4sfiw50QhgH4dSiW3+lNSN6VvajcXuIlaOTpGCNn3mjKh
+/t68nZq/g0u6/7zekKaWE0ipnLAd0zp1jhU1Fcfns5FZucw/X7rZhm3TME91uUus8Cz5sZ/MCTL
uDKDMYVwDfJVHM1XUX/kdfw68LfLlqY3HksYB0wEa3NEwMUaXGKXJE33txbKGzSYCi0jRfx2oIbw
OFNF7kSepvaiDk7VSbnrWJ4VJDfez5kFQtkW7FZKUQTcjDZto9HxD2bUlezsqyrna4XbiqA2j/0k
2W0xtGBU3v3DR41EZad+YdOmFEowH3gN2iQFa4M3/QRKsim/uSy7Mt1+DCbwmQ6dKsGxeAi9bsag
QlsLvOFn9Z1eQqsTyoqXyDZPPhDcOsiqW8h5tASJ87DaX8yjsnbv6sx/e0dhi5s1IWTAVmoDhNn3
uaqTFIqa0f2GvyJTlA6tllj0/bMKb5f9ahDz7LG19MBnVesFlXSYD6Al2E9HemuOFxr94Dcfi4/8
DT4o/hynXCWhrmlioYplIc4WlDUV0mi6oXVUT7ZvQUuFI5hO/ol7EHL5+jserCM6zpncAeom7Dng
86ROAvnCeneVDV8jguO84CcTf8fRb2keMjyopQ8F1bneVFYUAZZ+ATmrFrXCr+6FOCp2/d05grNq
9hYQHIdymq25DrqRglp3IO9Yyaq9r+A2gQZlycVhv+7TF8poB+fNHBAW3m5mUK2jBiKCCYYjhBvL
7fGtPfExgCuVgDhwgaupygFRm8tF7jVIam2U9g/e24+L6OXcTEoUqA9BuLivov/TRYeLYjHf15My
uXZ7ioNr4fLrIdB68X0GtZarNKF9fuwGhLmYRvQj8hCAwOysn36WyZ/8VLST9fDZQ8xr1VDJSISz
Nl+NPpSSJfvhEE5YtpVYz3XdS/XTSIyN3h76Q7UqH52oiAohoATlO7/JXy45p4ONoLsKert/qbh0
LB30CXhISTFv6jvOb+NPXtD5dxn4F7Kp8/nCTl9b/fq1d5WHMe1tT0UcSjc/5+W1IxB+oxYy+4ZF
gPDHD9oPRBMMcp+W/jCygIfpx7p6wNbOGqQy/+gtbu8tQIWJ06nj3EzrczMmaRLeUhIypCrRGzhq
MJdle5VrTvYKtqh564vB5HcQPbkcZGeVxYEEccHmfU+yGrxl1MFriOlKmx/tmXMwnBRZonxb5HEi
tMwHYmt27z21Nxk8HmQOAdZPd10rH/jdvOz+leSl3s74VQHrXjgoEJ6Ui00sBbfLM0LyUOn/s1Fb
f2iqUzidjmhFmodxxb8i9BXmExurutXfN8cbSNjYyE/9waru/fgtUAL/dmXBS2bVx1uHc1zyzRGs
u2lLhqyvWpF2ZSsZ4B73MfQO3dVAuuk0IkTaUghcyWSEVUbPPAE3Ps5QA4/z42S7koiPh8LNqvwK
ScVH3DftX2eqP1MGjtorwrHUzxTRX4Fs3r1KZ/qqpqdBQ0qQktJUGPBBmvDl+Gex5yaSdU3ix7KF
cgX3F7Zuj4EuZ9jHF6/2gU1u2KKCxwIjxQoxUwt8/P4GafGWT8gV4KZcKNMglHd1PIKfs0/SwRe/
lPTclZZc8QxDPJzCUHF+B0ykdvN3np0fgLyyk6dhN1k0YE3l9zA4rsVmGcrExBchV5fMLlpdzLuW
AyoPfaLdK5a7SDyJitkm5cWQlwoCvGK6eDa8Cr4sWst7N6B/QnmTZaQKk5eNzi2YzMMyHmwTK+PB
DCIDbmDaE/M1FkHOaVC7D2dLL/nc4esdvv8zwoGzTsdpe+h9Yx9QhNcZgkAcqcaT/qwof/9WhH9z
P570ag7qIEeztEKsplUpTRn9Q7hpsNfmx62J95uUqvaMc5mk+y3jXP1nlKxPteI4jEwn6zKFcht5
dudTGjsAtZOHnUBWJ7d0bNeDq8VC4un/uzs+ihICGvmDmxHVibOWRvJDrLysFu2NrQfYcBJx0Z+C
Y/jtXC0seKurHPPkiAz2FGR75FqcgrqEuf/a5e6X5bAl5CzQtyp7NTMBKrcwJVju8Qngo5GvY6TW
ExfEOgSj2u/dPjZq6iVUbXNN0m537xxNyRkn4aC935hK945coZgSQVggQo2ydGf/WI61potGH09s
COtl+MCghK2U/bdeRF3w2LTcj3Mhrf13WyQt96PdQj/JQ22p13yoNJWMu+N6Z3yP2o18ZnhrelRV
x2ZtByjmhkqSDpKaddWomSIJbfSgsgG5XDrreqrQmBTP0e2acyABCraX0rvt2Bd9mF4+vXdknB4+
qOOVrUFLW2Wc6BhzBgCqkyKZco//r78E6IS+77mrd2uin0Geo5p2CAMDe7a91c3Ep0xn/6x6Fa1G
OJejcde9YPBPNdhBEJKW5MdSfA20pSRHVA+qF9V5FQqmYsIC/nl4AMp7HMLTlHP0rY3L4dUi80y0
HiRm+JgBC6qPjWEcQlMHhaPEI6IMI9rC7PXTYQ4i4nsAIsCQjGLXt4HNkTj8TpoUGaSK2Pga0dHH
+0hMxoMxvWhRvbw0O9nJMjzsTzDYNV2QhYJHQQSiiTXsi5okmE0sAFtEefjBwmODGQmS917BBsQo
riTb0xKOanOCbsa4de21PB9XDYqKijMZDoDDMwPWbv/1xNfTEQ2JlXn639Lpz1jj3EAGYqSQ7xVM
zexCSME1wVZlfo5pkNeI8wc0XFN7VcylJwQw+ciyumanXQhM//Pe6jSBF0ILRrWZ1YZlxSsRmXwL
w6MqRsxgpOwhGys7AG26UKwIZmP4GBRyDnaIQvCSxBxMvjmnw2UIt9O0a5bKYifsbtyT5PRajhMO
eZd/KFlm6213QSsNstpIwFo0IGkeeFH3N9uAe5YNMt5GH6UATbHrn+Y/ofwXbUZ+sbjxnxDf1l+B
/sJWrgyulaaK1fWC7OxR+lXev/LxjiY406LD7aW3KCn2LGxDmOjosdTJWUoVV31Gvaq4DWPBci6n
r0F9/0wpLaVesMryrzXOlV63Lx53lzMQc+dD199r2HE9b1nPBCV/DG21k6/eRHem1DkOtXa71MzX
w4/K7rfWvq+Z6Y8X0qKKWhrO3A3Kjg/yTTT1o1v8UZ3IM5CHf2ydg6klK7wltWs86p8YrRBHDS93
zLC4pz0LJsXg29j8NuN+xd0ZnGWobDiVmIksJWvBwurwC30PWJN80OK4M8FL6l7UdfZ5BrzjSpdM
iHcgW/hOrWSkDAedjhltZthYQ9giOtg07UXh8z/KkzbHYt8rw7cLcFhxbccFUOdEZjfMxg3LwRWB
T1WzNw7ljiRayoEeq+JB3UFquITU8H3RYKIZNB62h+UeMSP01q6Zyb2JJvroMHyZ79WVKbPE1C8j
Y+ypWPsrzAQ+XrKc9rkyl8HXQAbKA5czY4il/IKPuUpEp5qUOcsJWnb6/sCGFePbsXU2nyM6uqQG
/GGPEeLUm8YMxlER0M0s/gmVc+QMusmt30w1EixtPZaxubJ12Z6YZtm2QpZpQGR+CSBbh05zN51q
USJQ2d3u0mEJexl1nYHbRLc7+e3lI0HUqrAuwynrUMlFJJHwDUveEPW0FtKeWjs8r0VrK51GFpwz
H0ONRXUj/2EpmmXJFP3knN8taAuhdRMFo1T1dFOIG+/CIj/oPUOo6qNLZZTNep1k/uDHs0olN9kf
FEMNjf5NQJ3t8gkQUnoWacP2ejRSr2Xoc61VD221a+i/KP2RNgIa1eLmrN8/epZ5oWCesmgt38iC
SwhG8cSQEbhm9iFP/BADxc19R/etNRPXtiMXeZK7nKQwm9/MLL45ZAZtic89rT278Ld1llg6B3ML
byH04Uenb94F9xQJtTAuegGBaIHg8CsnPM9Vu369lYNwR35J8zDCAv7htLgrYiMIE9TP5UoiFi6+
hRMpRl4Sg9X7Mqxkllh48bMgVqf3zp3VWBLa4BH354Kv6PZlspwFiqzFLFODYQxkZdlgDHxCi01r
QBwJ7dLP+iZpIOMRmFllU+O9N6kz0GZhi+jSd+VZKuSULuIJUrtkN1WtEuUFcMxzTzfRl9yIdjrM
OCC6ObIXG9HKuYIK2exRALvVwkBgxqOeHpqmed2xLQ2LRBYiz/YzVzUq8cI4y14y+5T1U6zpfrAe
SdTYx3VtqY4CAzuAXI0IRNZ57sSV6qwOd8RuD2Cwu2cZO0dP8/KHwWKMrXsO1Iok6Aaj76k4PVN4
wdCJ6wlc3pfvTBAb/Zkj8fguAqt1me9hK1PIYCm7IavsXqBPLHG2ZL+uUszJVJsWFWvumaeaVW1Y
FYZamD0NwQEBsiCgcd9WtUMkzZTbWFB0nzf31zm0Ir7NAw3cjbnWf8fG17qjPaxK0NMUEZhrx6rX
QYemiM/XqUjjGCV+czFXTDhEavpwai7fSkNHuTXTOR+WzQxBDZv9DUbHsCZUTnyRDshjfIxUYUc/
JQcM/8Kh1i+OTeBWFJa1GiBtcTxx336e2skdNZUqmcwbg0EVL1XjPE/8dQEEjBGgNlPwx+DzUE4p
1rIbbHgF5lFvSPh4P0ApZ2VpJiY93rzf9eX04z2UxLDZZQjOpQ4qODmCg0EdNfIastFLwlzB9Gu7
az07mleIlLKm0CRMGoeZAq5nWQ42VKd4l4+6DIqgw39QeYn6Ugq18mc1NU6Un6ro6hburv/LHXn+
ZkZsXi19I8vto2E+fzrPqNFxWgNJzkOGKwG+yd4lj55e7fhY22JGTdNQM6MOYlFrgU9iXfKOIhMU
zaJjuUeg0VCC6XbzYc/c8COK2Yd11Rro8h+8PJOINwp3WA+PZIkiLwt9izxnyU1RUPHpNvmu1w7o
OsQ6kDcD36EMgzmiRRP58rYxtgZtgvcRBpY2WSHuiT/3IUdQ/rgVoeCYekixrZpMqHkHKa0LA05S
vt3O9yGebCg247mUn6ambiGlSIVNxk9vk8ZHUnzGsPniiv4jycCZvW5GBVUdNeTXyl0ryKhtUK2y
JSA+56aMKFnBCWArLlz4uhNNBFIqFSoWZxxdM3nMq9wJEH46rV/luu7yyugoFI8QhcSy9sM90rju
kLuO7yv9GgflQ4Vpz8+Ou/5r+XrjSZ2eqWTZL0lgfmzHTDxJrBTAqesKvnqLGxIafduLBwEVqQiB
C91iZWvwoLpuwHlGC+qUJj5Ni0B0locdZ477p6JmWxn2vBdhywcx2E+c0TFFIwfHUgRymf/gqPkP
E5wc6eq5m8XaH4OH066k9QpO25iTvVYij0pz5pEcEg/FWy6oVw1h04rwp5ECPC4bQx49b/K1c1m1
mj9jrLa8wrzQorJRqe14w0eSSF8ex7njSAJcVO5uaDipigUZtrOGz8uGk+NgylNowrCwLUxfjjgJ
FRckRRNrNvey6bEmrbbYBJwT/EgYdjRxKfZBNjS4YjSzTjEgK52TcgTeuEqGjy8XqvE1ym/e8RNr
F0I9nH0J0/ijOG1LHgl8Riypq8zwxKcJzONY2Y1E7LUDG2lRPvmSXt9VOtzyl5JPXyNO976dUwp2
BmDxATJSZcB48/Eoc/7hAkFbzOcTzRgHr5W7/c238THlMpFu9KWA91/+Cno9uvOo8ZjCfc/gnXGD
Cnvh4tRz99jP0/cLXJw2+4rlvQYcU3RGxvI5Fb/wVtgzqw+u/ivp5X/Thj+0TsMyIMazxbM60Vhg
o9aXvCUZY4oUG0k7LGuK2vzmGeaPBxtqj2Se/19F7XRcPCmpRVvZWX3vopp7brgLma184Viv7WiB
7pR+86D0PfzMN0xGbstqu3BxpFZbxXHIMlJvo219vYGIiw7Huu0DIDUG8lCn45xlHYdpPvr2/tBv
eH5T4LDsu6wboksIpYgxW6ig0iLeni+MrXcftkG2x+0jY41++ZXP3QTwyDp0RA9Q8334lZocyWvD
ZaT1PJZ6PgNBfAN1JeujMxfbRA17Uxprv0Lyqre5W2V2UL4IAdBqmP+oly7pnYaEHwDwv8wqnkBA
Lgda/t/LSygBpBUR86IGtaMYLWRem3pejnUHS+6+JczdKiqa5vWGTw4RvgH07ku78h5J6G9+wSd/
Bv/eAFV8h17YWB1yTevq70FD32NLrSKRkZkZx9tWs+eLUWPDeeAttAKAonoUygFyWhChLM8JeHFa
u+MGt1L83dfgpuBbi98frmRYGlxr0yzu7iWf/5yhHObwk8V+Dpi+etIprKjCG9+/Gtom5X7e7ZR3
w/e/8S9XhRhq6ooKevQ9kN0dwZhtS6/EzhMyc6qcT3nNVy1eqsnc4NzOlAUrdxdfMbHqxVUgQHO2
+L6XZBfCO5REYQPuMMzBwAXcj+FERIGOqeSdaKYZSYLqTViDX3FTVyGW8O6ZDuTk0Llt9Qlh7gLK
wt7GOSpJ7TyeBv0u20VVDs+JguI4CML5wyHPltPzkGRsrbKqdEWJxUgCc07qu5sqH3BVrmQXpsFI
WORyuO6Gu3AYivbHedL544x+uh+4tPuBpbWMz+izXejaZBsd+UU5W8Ur6bVbBtQgL5jhEUja0f/c
S/6ql54WfZEROcRvlMhpkIRZe50CJkzZ1FKY8VL/VrnTGJqdBIkwuwHKMKBCgSvG45Vo6Olh0lwL
Q9QqGsNjgK2GjV2WoIk2nmCZALnxsj6MVkXx1fyrUjzO47kPEkZt+9nl34keCNfCrZ8hBoH9rexK
8SjLY2ObVLkmwxW78uUTicEVanNZCYdMAAugKTbDJnlc9E1IoKY1A/7xPBnBsFeJlZFC4bOvfc+j
flrhMaiNLJn3eFQrPSOGB/z3km5iPdzFl2xB2aeBOn6OasHLsCkqZozDAd36fb+8SrE6VGAJyljR
1jxVsZqJSsvzzttNLLAVqyoAXpk9AnK5G0+6Khz30xiqPvrzqs4cJRhcqnmZhvPVMq2SJC2vpINH
phINZaDTWgX7OoR02wTejvICSIoPAUzUUa11FqNQfrQhDuxxQaiZgEa7dPIP2nVdDkaYKfwH/0gB
lwn13aVyh2unSymi64lLYq1UDczi3Oz0UOaH1tQV5u6+xZtlFP/F1TY9HWvdmkDCBVPPXQnlw7yW
o59FdplaQqAcbNckVXddZt4QNdGPLgeWz38denlbc+kVKMW10YYMY8kxU0dZMLk+Uq9Sme/ly78S
/+RDGWd0xg28s3eB6PN5g8WyUlcqX7hH/IpPFGhmzfAq+CSwTuUK6jd6pR4CoNB4rGGPiBMzolOf
XBsPZFsk7z/T8Lu4msABM1Bbv/0gcElE4N/si2La6kakE/mW7zWaGNJ2JDaCMIpnr+dteiZNziFl
fqNRPJDYBOjHw7GnkTF1UpZRCNpZFXA401Zr3KJJkPipCzDkXksY9hgBbJMXJzo3sMBiOVDzuNG5
cj12OQIB/9pHz8iRVXJXmFkQAyA5utlo8aLbW09sDrH+n7AMdjiAotipisUT5KBDmueroKcoBw1K
rSUKfRzuShFKZv1sQfaPRdWU0wb01oXUp4XH+wi+jynL3AJgP+CukQD6REWd3bbviuHK8I2FixtJ
ONyzNZoMiSFULAAtoAJ4lJtct2+2Gp07pD5oeFBLZMa0TpLmIL8MstyjWZDtbwjrfpGtRVj7HqjV
x1BYfZcjp6Dxd2PLC+HjY2sKRWmC/hUpdrpNr96c/MVuYZOCeAbqnaPbDDDhUAFSdg4no/uJfLrq
36oiROnwuQk6svn5ru0oW7CIb7LBYuh7xA4b7nhdj2B+o0pZYigF07UgbXIrT36NX7dmYnGK1iR+
+9EEfXiQ/DbiemQohf95vn8lrvGwA8/pUL1XXopeYQyWkq/BxSbQm355YFleafn7PmJJ/hhILp7Q
iTk/ks0bhqRVOZ4BZecx5yt0jiieVFgaUHuWpZjkgqvqB3YaNh/2M3TpMJ+21tkJdVkZ2t5KZ/AO
39fHLQAIXcOasrij6bwwKuAvWpPiriZolVoFTpYKxnVZQQQb/rVFzoeW7tCapktYE6wAf26feDkn
GWz2cDYeCaSqxOODRuiWARIvSXo3YeAgdZgnPMveW/YsqEfarMtqdpWIHoU9YcDufJwKNXLzaaii
qZRaG2QzznsIREaPj3480+FbEJ9rTLXc1PCR+PJV6J38WlEuaS0S/ntgINbUOQdzbLvznmqujT8M
q4NxIgfW6CZp8KHpbINqoL8JFehtyivytFthnWSkVTPaD5EwLoEzuZatV2AHCrjpLA/Ae1Dt0Bui
Wl19SqXWjRFFBCVTKFcQ98LPhGNQphS+cBmQAV+tl87KtM482pZrfpuXkXZaUWPznKD4BZQxb3a4
hO78Oj8414cgEEcURtKtW8MDuzt4WOmujfmtYo0DKPS875E0T1RoS8tvpleWMhkycOF4xRhxnnlb
QtY8mxCr9C0bA7dJsE0EuwY6MmzZboXim4SmJtvQBIrQuZEbZVeaw3XKNUvV/hUAovOGSp2hp1Jr
A0K2Ji8rcgQBayYA2KKxeD0vhvgLLQHxJJwngoKDxfeXg1c4q48d5sYjiKrBo1zL0D7jxI1i0n78
2qD2vqCyepWZjhp48OaNfZOtKDsShIEFheVx7NYzHeeImkKSbwRXTemC7ybr0Hn/3JVc0k43D/Z6
CsdTM3Vn4ib79BKxif4/+jM9mIGP1ujZ4WFR7V9l2pw9/DP7PUzJEPQQXHBl2LdE/1uDONNgZJfj
+/P09vLt2uA2BdzEhkU9nauIqGc8kAXtQyQCBPVC75+SD8GXkFnM8fDinkusY0WChunwo11BMOpn
63Y9K/1U014VMETDksmaqjyDXag1esN9qbEM7inZ2cPm7k2rr7hVqsj/nCYE5GhRZ9uDrdpD3OrS
clqvF8kAx0OpNmBPI034HDfsKGeI2HQojTb+g+Jk4T9jFOr0JVGcwkqy1h7tA2J6alI76NG7ezFy
8r4JrFBwfIgKxUgv838Lo4xKX0kAilqwTqIn8VZjI9Wpxz8Ry4XsAGdlPNvWTGWr729Q+NefX+LP
0+HYfyuLfYuPWSbqTQu2NKbPzSqNe2vnrg6JLke92+5ijFeFgCmvbjI+SB8TvviT+9IsbADrBAxr
8GK3lWv257bxCJGBa5RsfQmkmkO9IYFwrC5/vEgJAMQcQ5azgEZthrWeNxhZHE07HS6pT9zlg8aZ
XqoSc8vnA/TVqDeuiwyWR0/+CsQsgiDj/Hf6Ke6e72fpn/8lL3yx7eguJWMT4EHdZshdeKjV35NL
Uac+NEfVdBrtcEP1d5NoCqzEHvnnQXbOxqdLiOws59o93NctMUt9dNGZm0SCQIMEXSxpykE9W/6Q
cyTx5W+6zabYE/x88LSvSl37gsc4tZOPCmqrV4nGBdiPYTfC7PveEASAL9BzBMj2xRvSVmuWMG+J
AaF/taoMojs+wmeRse8KXOOOaViTJFHwe48cVkekWVPVSFqgqv8PxdCHh4rcEuMG4MDBADyLW5WN
uzpBpT4zwnHPAMd4fqQ4OME83iFdtMJ0CPbhtHbx9yvavawcsrOO44cAveGzAmoa1NqH4azL4s4H
OqDy6X36oKv26tQXviuBTsyr5PWXU3vdC8WRb7b6yjg/3HvBnC7QR3jnGYm6tDffcU80+IZ+YqXz
6IbPo3pvV/uaENEs2JE4Sw21JZQt1VdQNdXGvL232fWI7EH1WFd3nJVLSo9orMvPzrzAgDBtTu5e
8uwS5eEs2dRYzRM+Kd2Pcuz2yk9qLRI0JucqEoh2iEgggGhz01yNtBcKy3tmmbv7NUM9DwXHjY8S
sefM7w5EvdOHzn9BYJpXgTtyG2gIJMEvkj0B+ZSRgEagG8GCGr2pROuUi0SF91Zabg38FhqsiXId
iPCdmRWDPCx43E3aFaQYh606PeO7WNGv+1oiaPY9QvnRo5nOCoirGyUyiBNaIASOlqMkxGy6TTlF
5mE0hh/qIJ86VwUv2Bmi3jHfiKHSRN7g3RGunV56KqnIAUzTns0gSV28rJrXTc5C3QzLodqfWge7
6Z9udzHTTd1qCEHvC97I0uIb0GT3LGNF0puj+ezpJy8n6tQcfb87Is/u7VsreU7AKTreDVKnjG74
ONveIBcC8a9b1Poggv20yYYoCWkksPHwTFhworAqOPRJymEVfOcbOcUonr0xK/gM6uwtPwUiPDpg
8Eah8oqRr/qSeb+3P76XE9a1T+xal1sbMBkDMSSv2YqqUHyVLJ59SzlqPOeOrWJrQ2NtAw4MEG47
MqvXwN5i+2e7mzDkchafDkSS2tnII3XXmAN/6/DB66O2U/TOP/Uxw5EGG/fHvHXZMnrkvAw18thU
XdUIwSs8ftAxKpFwAS3+m6wvMfBvC9+7+xzhpINdEdPEx3+4kP8WwrbW+WZrj2lSneZlLDOih74V
Hm5187ACUO8tkwZVAMo6HTupV//Tbg+jCPvPhTgxgPXwdyYZKkAfwAUlqmBUZuQRc7zNdNaNS5EL
VIOuB7re+xx28rnedoSiphLBupRdp9K+SAtLkgv/s9T2G5t1WYw4nDlVX22syFjTCZUUwO+HGCi0
X2SriGln4cjmy0IKO3lS8WDlJhVRhZxhsH6X/PWtOMKgdwphFkVWM3uzYLXrm3N3DsLD6g7oJS1H
Z6W1E1sG8xiLnY6sCZzFm3UALKkyD6sNUIhCJLm8qbBIV5e25kdXXh9AMY0V7dh2TbQSUovy+vCx
Qy+qBRBp8sErpki4nw+n1RwYWUBpZhQ1dm5aNsW+P87P/8RjBZ2Iczwe10ZF4UUE6KCI133qdBLY
+yc9S24tSm7OSsY3D3h1npNpXX1DsaHLPTos8dkYkWnA++vMAvf9GR+eqjmKMhw8l2rLP1Uad5Eg
CDNM+G0LiYBEl0lBjuEOyx4N6aPgQGntIZj7g6ERW52awIWEi4p5CCqNKVhFZHbnneJnOaXqj7kx
GZJUjuF5FdocYRQbY+IE/njzfWDQXj9JJsgMXsDf717kHg9q0lv3NU0iSoBuHbiYAaxt95lhgX1Q
rDUyAF6IkBwzLzTM6N9s7d93lAIE3qLBAjzXviiFCtZph7tbkwFivzK9HNNVjblsNPPIf71+XcjZ
d/NABFja7k8hD9FP7Od7bzZSM2GFMtXO7svveAKuDJ1oprvG9HPfvwAGurjVOO2ymqC/9jDW/iU0
Va5rfEX2Lsg/zHdFNOXRZNGh73FEy6R6G+dtLotMqPy7dthS2r8HusSlbXONq7QCR2tewnaHz+4N
cd2cGRou+X0QMpIM9JJsN/f5Gvl4WR6A6JEYaWGHPcMukxvqitgsSBlqof7K4exOieMc8+OaO19x
f+QLsWbfxnSnD0akXWjWWWErVnGjmyqIA1oqEOsDrWjLI/+oPm6ntmZCXdh/cllgyJKldiOsWTI1
b/dsg4wd7R3c/nkegRP5gV/ES/uVNbPKfD/HGOmNVqx2WfEQcK8CezF90lukN3Lpx5U1Wz4dUqOm
rBt864l7HYuOsXQ09D6ixTZzA5mOX86MnFInbNFx/62UfQbozSzYnWoS82brM0SpYWaYQJR0MpJQ
ZT6ijkpjNTFOS2qIuQOgdgpQ+GX0GqtxL1BNcpTYSv+06shahdxaUPii92LRXVb46YxOgMG7TvmV
1d2KYfKaH0Ynehi2CyH/VQibkJqNyfAZv7pQgbVUbB6BQagxaNu9c3xV2yamaGGk/u1cT4ErMYKM
3JCh7a/8NhY2//s+sGOp6WcS5hoUUYgV5eR2ChI3ham5IOPAGAYitB2xyMNyRkkEK6JznM+u25Gv
goY9DdluQ6Cv1/kuhk5XYhIhcFGnTwS/69vFyv0mwhI8lIYHL5Rip0fHoLG6N0/Oa6AAxXK3z23b
UIPQgJzfQman6aPNsVSoVxBl7SiJltayPhH/iA002XycdMGZGR5jzZPz/ZbTtGg5I8C8ZiTDaUjc
4m+iOIfQfd8dQdxMx+hjE3/z5EDMCGeP/dle7kR4czLOB3lWAsbixVCD7EcIaNWTisQy8O2Dk29v
xrsS3uJ5nhaL9SeIBl+1JzFIb0tz+wczA+CMU866LPMqJlVeR/n0dGhlV9MWaOwodmdhZ6r4D2EE
OQDbMIDlUsgtjsAzqkik3MwawHcBx5j2/zAmoy4bDELD9lhnPdneAEzmCw9NJUZ2mY5BXmjYPxMr
K2d8kky3vO9XaDz/OyCssFrVQ9AMF4eJVMfh8VNYTj2DHAebUCZPaF666FMQ1WBZinwp2KsVs0vP
tZ5oirOJV4mkBpHWd7jTP28Fumuc+rT+iFqJUtkdFISGPr7ycMb+dfKNIVrhp7vaKJtSz6G3qUp0
3m79e6HZWNRbZ5bKKktDgApNsY0xDLBK78eYiaxi4zxG6v0XE07TcvJwJIZl8Lz/TTpMJkz/8qJY
j18BmVAZpsdBp95MAhd58HnBL9u5YGhWYyksBL+fPoFFs4IRP6CFfgRJa4KFuuv33ZSENZyXAHWQ
0POnIK4zk6zO1xXLDjC/mhSNwQHiLO0b3myo2rOcBPJL/Fk1sebTK8WTPDNn0yCsjGeBZPGWDDNP
MYoNBo+CgQSNAvCOpOy4zcymh1QE8VkzJLqnv3QBU4ZBVI2wuvmIvCWVvWfK33QP8UBg+s5x6Okl
IPvzWvcgxHbFf9MCN/MTRXcXPePfZxQ/LGb+xCbGdK7PgqSO7hKzb95cMV2vH0qedTZaU9kiYIai
8c4HVYA/GbFbiNIXmcaSj6c0cO7R+y1kXEKC8vrR8DyO9KvFbZ+Ie/OmxkZa6OS/7mTJnn4Ppunz
uTJHwlJFE+Rd/nUbxXoDngpZ9PffnkG6rn59pZYUnqGp9kEjTauGPSaBrW74y+gmGIJy+b2KqK8h
4K/XVfssH9VHvzby2IJY810LHmZbiJbT3bMN83TajIuMhYcIii0L6CJ7+iDwctq8WZ2z8KPDLu3S
rA6twfVpUdkhbFwcVS35oxWG4VgSBQGArIRwvFZFZrGGW8FywQKwn86zddIfw4Y/hv7dYE6yxCG/
5GGaaN38sdIcppKuC5iEGJXyRHW3zCov+/N3RmYR3bAFDM1bP36i1CG+ze3ECwRJf6bD/SRZk2Nd
toFJo+ZtR+5Qf9lyKLUmqHXsTpC+d3hJ8vcmAGds5TrqpyaZKtJH/H4ItF+qwLMRdNO5re9wA+Qr
sASQZWv/y/sg2CwEJ0mS0NrbI95uoyO908SGlwn0sws0NlPB7nui9mNIaq0WPRnDIpYFXJqA4dA7
IoSy8wKydGWt0oes0AHVNyl+iV71G1kExWNBFziIVPErQga1Ksdci5ez6rjhlV/5LmQ3IdGaHLa4
2RAg4aQKmd1WmyKWBd2X0ZWXKChlKbg3l2jljsqzP88S6rtd4HrqD7kmsMVq01bY+PspTi9kWy+r
Fj6Qglz04QD5moF7VM//gqDHWbAlav55ez9F8RgcAfZ6wxlve9JWzdWobkBmLrdC20KeJhgfxO9K
KsBNypWQLDXgjIdRASad9rYNRB2nGmwUjui8ckKmtxPV48ZW1PpJsc5vhSaUh6ghQOjcusWJFnzD
pSLwtpk8Vx50vIGEc7P8YduVdoeeYwNoX/9p+Jl3B0vdxBekh4RRe2qWNY697kZC3JFpSz/7kVW/
XD4wZ8SoHvFC8E8bBS1S3+suYlTm1/zhqmtYOzHOQCg4a+7Zkx0tnUcwMzDcYTAJl/1TxRmE4xHx
KDBDh5GRrKO6eVnheEoVfxOVqnNsZ5gK+G+KT1nKH8ODYSXoYmxKOKYH0tKycsmdP5vHZlxtpKNG
3NRk3aeQhB3dVbZSN/wb2oqnqCKwovMnnSE31BrbNsBOjMa9eg9PFhayzfOM2Ccuf1IKRK27QE4C
ImwDYm8jhXuABsYSMfJFPwBvsb/aiCJLPxGCU1ZPsSu52Dissht/GhTnDVteBt9CY+wPt1Lx6vhu
cUq61X3KOSo7sCt9yB13N7TQ3Xt0RyOz5tT3vqzEhM8p6UGYKoEWeYKg+MG5YFtsBB2qHz7u9g5Q
DZJsdWg2e2BSynFISQ08aMNO+aOQyggGSLR2exL3ZKLVoOfWdF0z+fcgAUzyEwT607jkVJQiHR8x
1AXGYdPLRfBEgpV9n0nq+1h1VYlQVcZGNzUqbv3rawvMvWco1NiFWHOh9DCUAIbaiZFnlnLGP0/r
Pwt53FdSz/fFS3w6ln1Ulu3ZTkkVT7Xs+Yj2ztzgKeurLDfWdycPbqDmukaA1azZ5cS6eF22yNjn
BPtEGy3TUg1moB6r7XS/fNjla+0mUTC9+eL+9xkinA4YTT/I2AzTJIdmE5lzl7zakDGb3CPv0SOC
NJTKbBQsJo+/8EOAd5qzW7ZsujECI2Kowefr6AiwZBvD2J8MwY9q+ejxrNOdkWTjCSzBb3yQXAbQ
H8hmezJxo/q26zeZnb9i1giSK4Wmzryxo5pIiA0Hy3Qq3LGw5y5wsrpNicqjLo73wMO8x87tKvjR
VOu3UtaEfit4ndEhVpH/W+k6hbO3r6TPzWh4NDWOGc2/1Zw6X3ZCfN8yLY3gNumfJyLTbTe7kjub
JUlB3E1bpVVjZM3K6mxXXh/aQJ569gEYkSnLql0Uzh2Q4UCUqhJQdOb1GxzcfG/PanziLKJrmTSQ
xefQDmIUhc0cVVZ+ZPiStJcprK4E4tmkHTAxX69QpcjPUeZslm/IqSsNw6gau6CzNCGcZrqhWGFJ
ZRIdPlYPAmt9cspShQ2RP8qjQkVBJYbKA+oYp+4I5A8zNfcLYc9MRXjXFTkeFcjMO+7VZuwtHknS
WOyN1wKajDw08vU1eJYLlsoA3BgbdzXPjzXAaTIZp8Br5n/t7ONuaYjSzqrku0QCUQIvfXWPdb1c
4z0eZd8rF00Ls0h0P8UazOJLLhUihFDxwY9dKRfuyWGuR/nD4BKoD9DyuRKWZk3ON6hb1Z8xSTBd
l0YXJW7YGdR+/jeMdfyLCQS4rsfzhyyUwKkYi9euumI/3afe6MOPvNtsmTw0FQle6A/pGl8cQQrR
9bX3BXnZs0SePkJmllXGbN0a1rULS0ZyQxKio7fOSo3t8FBayBBFhpS0KbhmQWvey8u3SvqfYxbm
fyIJB/38NnzqyuihSONjQucLwJxqrJBQspqIlt4eLAr7NNtKcN81bAWQd0ZJ/kayLt18KtyzuM/o
BynlT6dghZDfdSXG6WllQ/4W9NW7NtrIRcyDzT/tM+AtpIsN7xAMxMJPbYRK3GOYHHMI+pk3vO7Y
ndSeBPrC8yAAypz2MFfzsAagdK8bV376bKg5niPOSWrO7VUqYLOWJ0f3nOHHwcl23Qu1T+ELG49O
mCwVbFAn3m9oGvci+B96IgKkIYUybgWezBSQkkydySVuui0jl6KL2b7p6VBdT0sudrBq074CUFqa
uZl0U12QcyV3xAdzyY+lvicB5Qkw6rpunNguctgDCJJdG0GpRmcJmG/y1OWrSWX4pKbbD+yN8Xx0
xu4IHeLsjF+xEc4Os5ME4PRmdOe8OXjBxZtOHUu0W3Oc58XCY3REuhBY0HeX9cS0a1umYZLBfGZc
XGo++m7IbnUvncd9wTUBLZRlcq5GDsEYsszMJBzVUbFX6wpjDZBTO/XaFOZ5XfWEZ6Kg/4Y5en5g
xJM7nTVPT9OtKeJt1w8gabQ3qYuox+044jIoT2Mix3qdGdDdCuGM9XCrNF+6c3MCIcVw+vdfPK9l
J3YhqnNrNQrN7KGOCpAranaaLR40rpwO4w1vmGZRPKAeXQPAM67zv5jMyN63MH1m7EC84xO8t5FX
Sg0KFFj7RA1fgBx7v7jigXgQHvrobw1QvGlcri5Co9TLuZ/a7bkokhBibyPMVEq0pKGLWSmKdewW
qEQxFD3/XZbIxKspFqcOTRRaHZdpMoY0vAwemRubP2k4FVayZy+vU3xS+L1o0WaHGrDuW8GWnUEG
ON+kH05sk0Yrro0HA2BPN0JqscsdCXLauB330vQBmPl9POo+sbJTbb5TGmIxRCExt6VAxVjuWBwy
TT9UfSFwdU2UoRTNtRoY92LpbsMpv/EHe6jNwF23mTSMeUBNi4f9VqzjCkYTSJTTT+GEO0FNXT0c
CV7kG5pb7Zf3UzNRfRpmYWStu4THRlxyoafNvzI5aoDIGBesB00lHOFOcXSL26+W5ld52z0sZ6xd
hWiUdxdsAGs/WVYQ5pxsSUQ5/alGzqCbekSY/GwrzPpIht7Fac2+dCLWndQqUjgwN4stKQ54xyW0
DabEpEVJiIyWSpwuqomWTbSGG/5cjyqaIqaTAh67PYG0dXKqtpnVp182+ZY2QzyQMTbNs4O0iGLx
abUOdgDxF76JkkNvmmfnwzO7V0hUYAGaJe6K/yeghzP21WwFC5Uyd+PZrW2ZflByUD5eKR3keu+R
OGEOESJHLhx/pK9nQYNMzUNe/BFFLtWfCMn12yXn4U4sdTIS3Pp2SGJfKDpT67GmFCOqG0YQ5Ahq
y3Hs4S5eAmdRBaIsCB+wOryF6xlONHAeimKAO1Hjoz1skbW2OLR5pG8xDGUj9UK98g2wDtrob0zE
Bq3jVbJuj9lxXd2M/89QRI0WxoS16LuZqI1HoR9tsyXuf0i6W7DWJziI/qUaxXdi3C4pHt6DLUP/
RyKyPFK9/IPz1zubq1wfNHpHhSIEF3uSzfg75gKoY2o0BlnqMjXUHCM4IEMDZSBpey55tptYEoUz
Zsk4WE4TopahMJ8fdoImagTgnBV1O5cxgmszksvsCQQ8a5aqPvPcFypS4tyD2c+C1TdmPpd9WgH0
rIt8SknO7uWfx66GePDSSSN+Kv+kCXGDDskDvO+L7OgxSYv4HCkWJzGJTHAji7shZ5pN1A5+YNSQ
OPlD+sZCHJ80uAP2mSF0Y4qKbHiaebwTxCVgVOUzjsQkOrdg50rhDzN3MTkVNrCn8lYy4jHf7IDD
3pa8DLj3iawxhMZwxa0qT/1dJFh7t2ih6WdQRA6bS2y6O262C6F+Z7HwYNhumqMeYIkLqEMQ4G3P
zNlbI0wB/fGALrEllUj2TTOkJmu5Yn4zvmwwYXF0cl6fO50z5pm2HiSHE257TLatebCY6yuJDKrx
gKVJNUAznKRpC+lSeb1PQvpPndGuWx6Pr3T/Ex9QUIm2cuwhdMJfozOWjbxM8Xo399vYvpkVz6KF
t77ypsdhKgb9eTN+Qx8kIAjFKVjLfQdSVCf3kYo8eyXY5nv4h+VVPVlaYYNIkLPXWkhSsdCAbGQ0
2PqB8XHiX7/Q1L7urL62fKxmzhiUGBoigvy3QQToYku/ZOI5YDWfdopJkxybFuGEjFN+pWk2Q/Nc
88/p7Ur7mocOuxdTXx+21DaOke6NqROdIYbxOkSDW/IXZnuYoACd372lr7AFGKN12hmDIJsRKg7R
/H8CtKaA1NhtyPGtwVdP9MFxKNmszWof9LZLflq+eL2EinsnZxUb5XTS+pNEKcer/ekae9BmKYmD
8/0023EryULyM/XoAezrbacDTGXKY7mlljL7Xq1qMeyv8+zTXSdWCf+T79actwrvzpY0kGJyvBCC
kOCjxVZUocKOpt3PGjHvTq0ikLE72ZAOaQTKx60NiMRT61HvbA+b+eXqzFzNNCiy7Mo5yJ2xSyn5
r98SRKvdBoBcKSLC65i46z5WGLE/vNlFg8WFf/H1daqMs2KJr5zPKbY1j8VTsE97tUyZeSC4OxJy
Flt3KBRPdh66YPPT2ONegm/abxVGpiw2wR4WPTnwP54ZM2fcjEMeOgAyrCx3lvAkZOdhGzoLVhFd
ewgCA6s15d9WlMkb96vHQJIl08cdP5Kvpnmqzx30IFc251hJ0K4PKF0+2hHbHk6h7Y0JEYisfgqn
SPQuB/kQY+kWvSJjB0/4sRa/qctuBwjvQI4Tjbqzejy4agUfkqszv3zF3QPuUX9RBViEZntUrjwT
mJJD6sCurEW3ln0wBQ3aG588wRlEF7KsNXWLn3/vU1+Y9wJty/5lMNwOdeA3TbJfeId3VX9nqWDU
1EdZbEyvyprnr6vfpX+JUKGEcaL16Oe0ZYD4twXB2K1pZam8MEXIBW6SJFhW0x4bL1wBC7jHD5N7
5I26h1Ts6LPHAL9Am26sZSnWMAw4ZhjhRPLjQvO3SzjSUdO/0Xp5CnB6LOoN7BirAB/xBpF3Yctj
IvHk+eIK9/jhLSVvNhWk8hdNq0KsrYKC2mjjIbeswNdksxeiRptaGgXq3bpcWklF8vPNT6waGZil
akhXlMd/i7C00DoBYSjjZhB5kRMpQJHAD2p9Xqfm7bNwwL0FEDYj5Q4uQnyPBjDQzmok5YzngUiM
rT7kqau1S6CfsTW8ySddfTNGiLK1C1hkAgvGBFkRXf/xkurX3jywuq0auLcsZ6cnb9Y1s+8XW9x+
6VFKs4L86ik4P/VorbFi9dn33/O0gKkFwBNtVetjP/9rW1jkXci6mOOx8t7T2/OsYdmYMQYUDaZq
VBGYdFxrtAY7ItmUrmPlU6jjNNJbbKvyyvQzePDimk0yOTZTmBQoT6mi58sR9NAMpI9OheLSY8Ff
8dDNYvO49EHkVR4Ipnjo3JbpOxvcNOjMYXPL9H2LqId/P2rnZMPzzqMeh4VCaGY1DvV+/5nsJiIN
c1M39My0QqBMKM68r5U6kdsoNkNjba30tSEhhbL7qAeIWyFzQ5nZr8vZ4HmgkhHK/RckCP7Ha0P2
Wxh++TT8b/6EdX/tHvUke4apXwd71/baY+o+Y5kFZabrZPaD7bEpDOL9paaKSVdScqr+GVEY4L5p
+awUDr6N3Xa4n1wzoIHYKh6YYKdVfMhwE1aOYr0x7VkshR9qFy1o+oXTUMrSFfJMMh4qHglhAk0j
Pmvjsh+O3z3HU7ewlMG4xubgNv5mwqPhv+RUiX8bqao8PtKE4YscEUT1hT2Ul85otxfN33jjqXd9
W1ZTee2SFp7/yi+7Pk9Vr6rpDGr+BCNDFL6hmgOLPf2XwbK9ZeF69UVgUKK3SZU8mFp8ofSmXb7q
DDNFdvkulqAL/OSD625/LYgJf3vmviiuf97PindcNwJRdWjqWzPE0BawUOLKp458LjHpvJm0OQ5Y
Vq4NBeydgcGJ1hB63kMUKr+piHym23VMrTlPLOdM7FC2b1jBk/rNhGjpL1WRSNSEecuPLbAg4djg
/0Zx1caxVJq3yiH8eoGy+ceSQzR2j/vw2DD/N0uBJdR9VIpzZnXbuDVepBQv6inocQDd/RV/afav
cn3uv8Nbbnoo4eEHIvc6re2pfcbAeY0fuRyUyJQMDsIyFgCzTxov/j9Vjigwb2ZfHbIrsWLFR5rQ
HX1wBdKS+6sZZ2JejGXtXlVsXEciJFteumLDiOJPo3wDjLpQGFNF4ST/mCmc2jQvPP1NR5wVMZ9c
9/+yV+huNtHjKBiMAX0nPxhIBjO+XDmfe0p7qhKimMgZ08ITgcMtneb5Bn8dooFZPDP0r+cqS08d
XkAjS+bh0jpN45TqaFNAnRVqHCginoIHARvap31ZgS5+aj3TMKsvvZzUB6PqfZGe8ODYlPjM1+Mh
qnVUGL7GIO0xDle+V+YTzYoZNN/Tv7IueQiPiGqyuEvr4yQ2zeaPWl10F2AfKiykNxNGRRz36O6F
WhqFBX6HLS3qlfpHjjb0Q9yzHQuXcXQ+Po4G6nnfrRKk3UBML18wBheO6y1cZCfpCdZGP7xOpLRV
8AdqZ1c500KgE0RA7v5+QT8AP3ZU992Ui0QgaaZ2xvw0P85UmP4wg3TfuIDoN4qOtLr05DRdelyg
CwZZ3FKFS5qSpXRSnvRYod68QbAB1qwDCTTC2R0g88LQJ2TP+VCYeSBZUDE4b0o1qjooBWw1HsdH
vaRxpF8Jfd43/yo+CoQg4ORLBIeqrYpSEvjSIElrFoeSTIj6dSZxaHVOgWdUgIjcP5itbR4mApXc
maez57deXBvmxvaJhB/djWRRkWvTif+pEHifDYkaBl/lG84ky7i8UmmmmYDIRKnFINSvQb+rJaIq
zW6HoCy9MdqdOZz14BYL1R5PFuYNP23s4AKgkvpMSRRILJm3tSd+R9P0RfAIDE53Omk00Mob1Fip
K3dINebNXaOf6fEJCmqoOVNZXOdKJns7yOaAUi8JFOiUSP+IJNjTnrLk/mvHnHsf9DKdDNXLlxM2
WrWiupGQi7gHA+4AtMYWBOv1WGvGxf2VXE3tHHVfv2DbFPhXpN//4DGbTk9Z5nv5hlKruffd4KrD
1YxY3a/lL6dTqiA+6xhAi3XHAvofmypL7bIPrrEQgxJmQPbF7AVwVl8gMSNz9pJ3R5aqCJ0Pxx5d
sLRpXp/QtFEoblO1hZvZO3YNB+S/ws1lpa8AYLIe4S5IjdFP/m9b6QdogP8ihXIwS6b19L6WrsVn
vTqW5Vj0BQDWJNIBpXLBoO8rcDGJS2WmqMzGjGt3mUClpAhIvg9JBJGHbtp0t5bFhHdcnyC8CeLj
Nr7NUY8bMDlZMduvm6MxfvE4zsMwA4t5PHyiuH5rAZAOpJ9YhoBThaS+oxKiQzmFzZh2NM+6tJ0h
8ei7S+AevOIF4LErcnQiyIK5mUeU+RBSBik5NTFZHszAshmlnNBFHlfFTrRVAMvlpj+J1wjP2Msx
kjoqJNr6QdqSicYj+wS15++2uVWf8YKfg3jbLy94Cz5q52PAUdZbR+9fyWRQ4r+YhjJ3tma1t/0l
U2lAyfmZvNtKGRcE7J3eAJm1wSAFtdufiA8Oh6V4MpKMqj4BTQo7rFT9ap4Ajn5pWNXCC/qJy3pc
aQefzmVK/vHEJmv2v5AZDiQ2x3Df2BHrLKg46V+z251fQbzgpX5v/THHPUyKWGGdbORlCj3A1ZO9
242CliCVT7McyL1AR9OfVHNXlQypA5dYn0Z3609luaG5jgJDu2d9sUoPMrc+Q76wiRRFAczwn1Bo
YroxtLdDSCpR/KtAa3ndDqM8fV/4cHBooak5hHJ5JFVqikKqJexR8MnBcySLJZu1fa4j840oS2OZ
l5HvmcbK26roFvfDvVEC3HO5aShpxsrttdpClxRyvmN1b6xpfAOMNNzlTfPZ7xSAi/PJF3Zj2a46
TJRM97GAsnjiipImfaAE+i8u8v/GfVRDWryH8tE+BPxm+WsuCypC7R74fdIfonEMoRkx5OBD9Ir3
nelsX1r5Iz+1pPCVjta9TY5upx3ZlIfrcxIttURrwam8GDMAj2inVUQrcvetY1jZIXeVKX7f4sZI
UPCQHEngiAhZvUXirj4roAFod4DX9hEAMHw1VrqSXAOb5GBTeHmlWQUnsPtlKj02aPjoJsK4Af14
296JgenYdGvWyJLGUQe4ah1ERL/sw0cAMN+Yogyc6OwX6Acs4Un2GlfciY/+aQpznMRIj9uFq4T1
ag5b8HzWtrIpJE0mOdTz18IyLAXCpRF1CuXMt7WlRnIMetB5rH/wRDD/ARHGT3tjiB0j4TBSzxfG
FYyOjlggnbihMwnew8Ew+NWfSZWfgKF4CTAAevKtxbgwI8rmNoajcMp4l6x1sI5j28SMMaBS94u/
28egjdsBf7WJhd2bZ5feqvmYiiDKQOM8iMa9zyOxxy1ngyLSte6Hd9DDVG6asqj5j27E88SDCnxW
RYYe+qp/WlfTJlK7A8l0hdRCRlmWj0d2SQDksPLjLmvgBCQ0md/KSD4UiotmOqJQycbTxnyKsKNq
DVf0bAZ9cN6SG4OJpYLZ9J3UO4SaF57S+/oFgXCTpqo+rdF/IFTSXjdHWCI3E70C73gqH3KUg7Y7
GJZ621JOfFgvHSQXK/jfmrb5ritr/183Jb017r/Y3HY2txoopOF6R5V/k/0RCbXTjSizPzdhOQw7
Uoy6uIdt3eDsHI9AUE4au7/+xS6dJ9sMm2F2RBqckbPZrvp8C8Ie6fpA/2X5tc3SRj0Ra/A9lfJF
fUWbfkXlCMDia/F4hTxqWDDU/cpTuraSivmF4b2TYj+WF/9eilDq5fMYduJKOhZZKebLbTczKz+X
ptbS/1q5QH2wiMvcx8pKdGDarH3M1TnM01j9wPMFJ1BmgrPHZybbStdLuNsRDzjVSpXfjpJdfdJb
uU+k7nA3hK1r27DItTlXywifMMEkVggH6p4zkA+FOiRaVjBDaba68MPxFqV3GmdGZMn93ex2E61q
DOW/9hbTs6jATTnHCkbA9pAeYUrLtctG0Nxk6iiEPCwzu4QgUm3gFw0uuNhfNtpAbVYCL/OKZ18+
ArUAH5EthMxmYNWYKm9ftKdMRH7bqjEtc6QAkPWHZZdjYXqYXIcfJQqWIz4t4Qil8CfyXfSCfCsl
Wqzbo69Gyw1gD8fAfGy13NHLNttUlkpwFTC2Hk1+jfkpckIOnhsa7ep6Oj45vQsX8bsh8FCdTOeu
O1SNNFKowyEAoG9owxka6yDLVngIjMtxtsEgnc2O11MLx4r2Iwg46z60pESRaIAo88iG8fJMFAAK
WdbPO1CySaRpRWHAWc2DDPHwYWpdhC5GPm/sPFnaQYtsga9HU5elcncG7LrBVK5raq+nJ13inYaR
mu39uy9/IJ+UdcpRA8knZuJq1/Z+0UYXwTVKpzlJne7wnYeZGEWcBAHF8Z9376jHPuyHk3qFRzuh
fEvIAn7JPZGQjfYOnzDJr2Dr9FGGPrgz7/dLtrBDPKBSlndyXJHWnamqBdFsnNxGMov7GkJbHSi9
+ar6mBMli50di8tuJfd9r2a/nuwfob4BxZIiY7oHmeA5UJV3fF725bdm7BTi78lWj2jchB+YYPSq
ORL8LgixOiCL+z52T6btykXB24BY/O69XonIlfVGu+S5RhIAlfhp1f8TiUFD0foLKlbV0QJpUar2
mkSWZLoVgmecHAGDFNFnVlmpSq9eUq+EKnndIBmPIbLwwivzy1cQxPhVSn/dDeovoIPCmLzaocw8
bufy5nKJihA8jNlFYmltmENmKsxlcgMo58FoYkOvBD8ePXCsTK282q608YEdbhFeuPXXKRH3mkzq
ZiMhwZAICvUHevkJJGvFG1rQe2+yq2y1zuARc9ox9cImKjdmFKwxHWHKdnHoaMl0kmEQFNB4Z3YM
JLnx8cOTu13rjwhvDU868x7hXtA7/k51ObfuhBGHFwSOqn3VSakbm0jGSUtgqsHJZtnDJ1yMHKJ8
kcvhI9J0p1OY2jaoe6+snln6OAk6dKZbx9PHq3xTUCHt2bcrQA2UwcHDN7L//quZ7bIQICePsEwj
RK8qFA5dhsVaLMD+EV5pg1B1KaresPtXUtYSxzhCDaTKxaui1Of25FfYUHgb19PzPQ+RO8VP0l7q
KcKCOys4jbev1piexlwmtyF/oaYAQqPEr5ySZU+4axopaR+HoFxj4D/ZYjH00/lPWVQuKB17+up0
34ZAD0ry7S3zJBgvORSXc3STr3TiriivL1uk9HdtvbykofL8GNd/a57c/UPBZJdldKSbf/B2V93v
zAUpsW5cUab11rgBbZOdsFTeCGAm/z3A2xtXRjz3U/rRpwEAwvUu62kVLZZ7/J+yLxD77gDqBYJf
lVrEBm+gmlIX7JHZiVerCYjiH23JhCbfNkPc0mfJdYpVw9dTwVxe4/0a5uopzA8/ECaBErz2Abse
TyaXeCnZmSDB+U0CGUS9ZDEyG70ARrTzhLzUAI0vAFNAnCcXknqaS8LhBENgd4ryyYOF2fbZS/0R
kA9g0Khp8Zh0gvt1358mDPXWphCd5U2YICFICTVDnHdeIajDLYH1pwK4QaY6yJOkuCaWyncJmJV8
CgdOG8J5hC3P3BIGc9YtytS4X8LtfuHJO728JKQbYwLb+ZctiyxK+afv66N2nHdj1wBKJWBY7Ov/
buZvfYGHThdppW6sXhH9Pq8+0MDdc9qEhroMNX/fbhGEabJrRaM+h0uk4N8qap7MAgeje++0nGhi
S4Jk7fGvb+yPalLB7OGi4O12P7rpIjUf6bmMfr5fJrUunl32ug6MWyDYfQsgz1YhTM+69RTFjwwK
hiGVGB+OYawuFGleYnCPS482PBFDYzWyI2Z9+2XDKQCXMVmgWygiqwUZOQV18KJUIBeanPnAbrMT
LyV5XUNb7V+RW8Q0XL0DGMFOAsx7o9vt7HkX4ccqaKpQgttbv7jTH3GC66n0tFtEcMbarqvfEnyO
+gB7lBRN7sPF6ljt/K7ltVPeN4+uBmrRzmX6KFuUKX8RDB5h8CxBeCfAJIKseGgtP0JPFMjCWNFK
x5yp6BDJMONjxZfXJDu3Yoop8YWgUzRVOQDXnX5/p6lNcnk9KQaZxifUUt0cDUSWRTNXdLJJDYIF
R0/+blGq/L82DuLeMhnjzvBcZkIZNRjp8DuKpqznZF5AENDY3fYmRzozq3V+wm1WLyOuNEw3lgIT
x5bhlj5BV+/WgMYLFXH/Gg30ZhG77/Wvqy9ECnWTuu2y9n7dzAtTyM88vy8HgSRJl9KUrD4xstSN
olL88PT72xmKOi1wbNfzXGcqBxoA2ClIo3SmbzgOX97eJha4iAOqMYoCt6qTGVGmL3i+OzhYyhtE
3qdBQk+MFgfURQJg6uxCqMYVMw8YK5+EevITjzgfvaftF9fVKMoOBmFpFiCtSQ3wm2qUpG0qxg+k
VbwRNo1Esut3OC4vZxOcBs0pWtsxR1ueX5NSa/XcJtlo4Y2fgO8f6nN+9mBsgH5rCOS6mUyeaaOV
dVrEKb/7q0qB/M7UsgpRDEm08yngcM3N4qB7S5uFmN0vjuyUT3tZtjCDcxKU7RY8HqSpGHwFcLH6
MVF/9nUlGE2AeyvjAYH6chHr+AaQcgLpdFe6QwyNth+ZL5fCWRPxXFx/6e1OzVxcDa1QI9N0OF/w
WPH0nd/Y/Hv66gJkPdCLU5Ogh49J+jFAMvvd7g3E7UdYWbMAbtFp5+Vz1Ln6NQpD3MRKjv9RpACB
CEzCqr1xcVmEVsz3GCuGVjqxGhxLTJvGGYDb161hdypVBmW5gHJKAHdxrQaFfTEXxkSgMfD2KkSd
zihCtm8fo9H+jBkkZCYHbFdZZdm3qt7iLlISLDxOwvin6I+0MFdiHvgeJl3ujEx4Eup3OqCVk+za
fBQZ0eKiVO/yTV3RkPpWwF0m6KyWyq5VInMqs0rXWHUMN+ZPY47fwfoEfhRZ8xbv8muJ2rQq8m0g
gGCFmE+NawZD8MqHq2rcNro8XtWwoDkwFZ5FAz67I9KJXMDqqPTqcbKPMJjYgOXUlSLNe7kgBaZo
E80y9BrudQzuBEfTQPKlJLXuEdorWqPQiUUpeSb5koI1EgDCiBq7lJ2Y/Jh4VnOjXiesUnPHrIYa
SEJYkWSls6yir6aRc/lSSDY8JRCbasaA2w0727kdxbu74Sy1edj4vArF1z6M/QK3FWgRuIF+WC9Q
FFOBGQ3cL6uyuSoxXBO6QfQpNwzz2+Rc4LbXXR7aymdK8SrZ/XI1esuSQUndbQ/OyN710bukZNdR
E6ttZ/pKFc9Loogbj1qKBa2VIYickHFeGoNKpTyTTqoCNS4r2c02atEZmzRPU//bbXHKh5p6prEs
U3Qh2dIM5blvBK2/KfdWeGWh4w1QNAK8HVd3+zU5q+vBP/XIkHbuW/qRoWgBYmQZu7dVAMYSGED/
Eftke22Zs8nXDBY6lwsPUgMuHGS2X7Q6GutTyjy5/DzTnEqfeTI6/GfOpGL7hTXlzNgaQ/xNtHzj
yZ9NJ4YfnmjYOPWpP9ayQRBhhMSF/67mxaH+xVKW/+S7JqKJsL9MDkYfaxntKgNLCy5ZIrF3A790
795Leev2eEVnUcfSmkRe8rBsNihpxeco9RRhuLf+i5EvIXDO0BaHxYI8sRRXoeJsxeoafK3BMokG
BoKTpbwyP66wBfKQ4OSSl+rHNQSaVeF/xuodwgfsPA5ofknsDh40DEJwvvy5ju5/LjyZGx6p2NXf
xKFZr89MO1uJbxt9Jzv9fEzlNpx2APNTHzOipfeLCbUvez1R38LPb6L6Dkt2ZgZ7kRkgvzg3/T1o
0I6IgbzY3iHktxgiUTH+sPLCTlavZKwQ8+o+FQMODQn3TTwhJNYkHrEXp1zmJLe32xHwPmJ5rn8J
+t8BRXKhl3dSme+/QwiGmJgNyUWIcD+KfvSJEN2O4pcT2I65y2pTr9W40jzOKb8AGyYaGVWwo0YT
Q5GjVX98dBkRwdPiapE95g5fILdWbGcHMoQmT8MXlMa+ipaPpYbwF0FMyYfq0SzzQMxI3FH/6MlD
jl76cqiwfdCPm/EwVkDf/6aRZxJkggyBlBdlCiDjgTRFu4hc+HP0x4Evmj9dAs23bAI9eLbhZ+fC
1RzPNrYtVSZIw1mc4cWdC4TIwLo4FsS3VinmpSQznKTE7dx4OsQO/+zXfBmA623RVTPW4kThPJch
Vbo6h/T8vPV4E2DVoq1qBalGlESPB4Jzkc85HCr9ZoSahJiitP8Zv9z+xDtqXBvb+D5Z8hC4HCm9
sQ561P7e+jZmuLBVLJSo34xOGvnupAxbz4AD49aMBdk2UeW1lzBLk0tO24b0/hu1jduQexULapK5
hb5Y2rnHpOCzZL8UTraE8Ip8XFUcG4X6DRCRDDKYF5c5sMDETJS8/ROj8MXYbQl1GXAgqqZxcLC/
QruPv/3EjMiSXEMS2F5/CE0SLSXcL22kpVwf6qBXvn1lILDNPRS5dHlpgLkKz8R1ggzxdgXNNk12
6wBpwqkyvXDxC01qpm4Vkh4mbxr0B+4il2W1HplFIif3Tv6doRvpO5Js8dVu0PqJuO1HHD3HFlBT
S57stt5Wo/X6DVbTpigy6pKyfkShWnkkpnVyOwXDqNM0b4EI6GSaiRdMaNTUFDFaWlRsRGO4a2zw
hNIHWFBskb9PNmnB7F0ew7AvfJ9iOwb5FgtEo1gExbOS3NI1+RewEpSbdYLIDXwgeJiO3QUOgEQS
9jdcUcfgCw39hhHAgGAbkNq8kbumxLOEqXGMD50VJalLszcRRc8bTpA6FoUguN/VbYZ+rN5j9j5/
5232fOOomeE31YcbKKIvRnsZNT2+LrI1/eO+3e66Vfig4SP1Vmlx4iNaB8ItUGhPXnrjEbbxF8JQ
J/SGi+X2vCTRFQXiVBEc6q/WUuYiqT7dTlW8idW48SW49yoTKpPoJKFlL/WcOTuSUOJTNYKLZ24I
WZlks5oLiwGU05g+QXirViVbBv8J9bIJcynOo3wJ5cq0y25uohj8Iwo67yl2GwC6kHqTatyam6IW
7PlmU8jeMl6QCD01O5IEHsadaWQeTIjjFhd3w/e4rLaSB19NWhywqh0wHM2QtDFaSJzEXGJADYEV
KEKQly0b/hLuybxdI7Mo/0CwOfPhCPUbDs1C4Hw1iENZpj8p6HH+VW27Mf0JWoHF97RWcj/KQEAl
jT23y/vWmVEPtn58PXXcYkKiWr9TV9OqI/+qNHM+OVjCifQzBpt1I3gwE+XltaelwBclJFFlOtFN
kjxOSoMPSj6gIOsyhN0Q6TYvmV8w7g7fWMrCpaXr9M+RFlmGhg2EAqYh/OzJ5Buwb+TuvWjKzvPM
tYzvPbr+CsVtRBCbRHoyXspYZQdLl1cLeZ0tTTrdw92DmAU4ikuSu7P4HkihCLJUP3GmmaRtc7t8
8eX6ACBnLJZHa0mLbqo+HOPIobEK22pSBRDme793oeTohS3WjfhanTL0Y1TakM74rd1frDt9Bpxa
3TFxfqNRSI6bTsX4vgZBVT+9nxSHfCzj2W9bL79apYhGi3dF2wTODc+/3bTzC1/wJ829nbnWyskf
+B7BVBthj1bUL/kvCXFRXkzZxdwv6k1Ab1DsTpte9iNasI/pVhaxbfswib0uQOgprQeZuZL+MqnN
UJ+HP5in3IPh7ObUDuVcjUAjUub/VKk+n4AbThDA8Ppkuubng3hovK7WQeGcVgV+jQMjq9zMXAPT
ChdXBz7b/g8z2ozXjHdgXOvKDremrthoGSnmWjmqcCciACgNXJ0mTXUz8GdW20lkwXP7WdOUdvn7
UG2mRES0FTnWTYRjEED/qSa2d/TomBNo9Acg6Zd/gDICNgR5IBJ8LWUc8R+stMMoPKlOvxRSasj5
FAKj8z+8fGc4H6PZ2GM3fwVnDgcYF5z9Vxb4d7btuLjo3kzgPkFsV3HtY+ww/Qc4/j80v+Irt/Id
FJdJRuVpMNyHconRGuTHRQMPNZd7Xw9J5VIOlaQOamD88bYRIryXy2il/5AHkKYFb/UHISqeyKPP
U5fKeDGENd6/TdE1qw8TszGph4BKhDKNgpBLfo28S+2Vn+XUe8y6xS1f1uQ7dkHafwCuAJPaX6Ib
pAKC5JgdwNk4qS770fl3wHsFaUjoBCVUkZYOM/MQKVre6vRzNul3p/TVm138RKhzAaqVUDb+b9s8
qXxs2AO6VdzQVbZ/BIcCPYh7kQoVwtbVQBOEbWJlCXUKflzOKajXnilfnxMjoUCygbOX3cn7evlk
kCTFI8iLgj+EaZL+rDrK0Ozi+nPLcJFrQDnkG+NgY57Je9xJMNHqALdrYH57YTQW3L8Yw7E2Q53m
RsL5X+fZYNMQLkdMcAQPYpvZRDDuLFv+Glt5ZkXOaFs4tOIbUFbfaIgXc4eanCzZnNkuPX3/+uMa
jQS27A61cRx3s9Y3q7kbngFmsF9ORFWIeiqVWE4quqXH1qMLvrtKa3D1m8t7Dca5cMhm/LCuOSez
rRswwW6lgfq+CTFJkyGy1GVSt+8KN6IYns/hG0esaXvUzfEpC/t8q8Jl7NQXLCdLbNNRV2nEmRNR
cGgEJhcl9k3JRMqa+0IFD8CFT+pnBUofDFQkJzdKmBunyIhvCE318f1noIHGuKpc/nNKy9sZYR5n
hSe9u+s0y4g/jggNvL78r43WXoytZoBPMQIDQmfFqakSUda+RBAgCzSjX+ZLKuQYVCOxRRUWSx6t
7LiceK3NJb7o/q+spda6/V32taquYnjoDFeiGAAYZgGM5/jdh8QHE0nYLhYv+w8ykAacnPBSgcS1
BwCQgEZqbzWLAki9LPFKFEgCV+FOGRS43VMW76u2sRvtw97/ifVNF0xxtHuI3ZFGbrh6dpAEuvBJ
stflbc8Y+bo1p4gAdfvMW/8wfsjMvDrr01O+vTq+1jHTJkFvfPZY/AV3DROQMG8Q9tKCaOjqUYtg
gTrHwUoTrZeWIh98Iwika5ZvS+jwzwQJO47IUrLMaLk6O/Kx5tVALiUPJAdsXT7owPFPObbLl1mY
eJtPxV3ZeRgu3YXtSIs6VkNLEbkQdAvGo6aoavDJyah3PuwvsiQGDOf0wuWiwvi5sOU0PSpbEmfW
Kih2b7cos6niBeFokSijuhCP2q5UIRPfQDWML1GfxDWWRCQVue6geW2aA8UxkpkQzaUEaouZ9nIu
IdCEIqjWTxSRzJEq+bnVntKkJAhxNlXHd8N23ke1TxcuZMUxx6DH1bEqCcxphf9B+cZYwKIMZaKI
lb1QrMm4V7f6i2j5bs5c503FCN4tim67SnRVSUzttIWzAJlyICvdE2jq7JGKT36nU7yDTDwkB6rr
BZ6b1MaUXLPFsgVuyUhx8S95He2OYsCHmR3V1X9yreXdAxunQsmhAXp9VV6AoegI8iCwroCMfPMD
UBIWLal2rkNi1Tz4qb2sgB8qDmzmrCR6Nd/eRmzwxCka4tiDjwswpUNsBS8/taQ2TitdRO80I8LY
AUzAlvwRjstbGHq5H4nX/WiXWVPBQVIbX24cRjvFFAs2T17kvmWPYP1ssv/lDK8pTpqgGgb3fzyA
aP7BwUkbsx5HVTCGDvyuKkxbVFYpXzTklVqk61f2Bq2fhbVHFTZhGc6gXLQZzA2HbXxvCOx+tXOz
B++ZPki/548DxeKRx85/o9zELTKWdyNbQgJA8Jcqx439tdgX3gdumdTNLmbFlWzJph7csufwZ/zX
3XkHtkns5ERpYj261RHPbR1VfQGWzTDX9GY2cBvx8QTlQJl68cbVV9PT1Wgifw/YVulbILiOPQU6
1ru+VQkCZETD9HsaGi81QZenLDD4aUI8R3MqQx3MSgpoiCw5vQfE6HN5EUq2s6SqAQF6yJhfRjVm
P1UZAk9tDr4ihjOJxjotV6HMcnnSWJDly6Y3OB8UWlxD7cwF8S5XGLxb2pLVqnqffLprCKt3Ny/A
pzSkVlJGW6RLdhMtbiimgQQXfyE56Fja2qf9Ffvw3tsCu2nl7FzVoq+YCC3Oi2A/zqFtUt0MyqOp
FbtQDNd1dycRIBxq+bIxSebRMYvwN5p2T3cIMIPKe09e9pcfB8ZUjv8bthZms+akrRXb/2HauKIU
l6nmwP6lhJoJy1Gr6sLtiO0+BEgRTiIHMTufaaRwPhQWWzs8wqCVjoD/Q4QHcUkW1j6IGMkQ+rZQ
oL3dw7GQXVRJIl82VlpE4SrGgHz+nqW7IhBGPnaDJ72LMkZygYprhnMM3YZGoO4Gla9FSIHemhxI
1GyeIq4ihJm0/bp1/XD+KaJ1j8TYkF5KlirKOPCyOwCOA2KKXjQhSgEbGcB4u2XfW+QHbBJt1UsQ
xkIMlB4G4L7PGISyv+AMTg4E44CgBTW8NmtDT9KrsB9v9cLb77vmxWDGOtGFIv5PuYuJ6b8Bun0B
LqOwMB5i3/ehKGxKB6N4AoS5dQ4ZKffqSab1Wq7iMLW+CNVZ2p2ceMZ43ZwndcVussTRZp66fFh7
Z4GnUmie+4YXIHMZGqhC+mQsq4h/3BlDSqm/KVMsvBHD75suuO12Cpj9GWWFLdtm67ZVKXz9rL0z
6KSZSCpBklmwI5IwsUA0Zu487OgMpDh/JdOqM2F8VRmDuJYGNZOqFFSqo7dyEGaDIJT547tDzTEd
2rIcmkZo7sTG03m6C31jvhB/A87HGStuo2IPaKrS4WNWMtU4XBv1WbY4+Sh6sU84ipObbgAQ97c8
JLka1Djhy18sos2AXTnP6qOyI48otK8TqgM14M7wpjvHL8xU7bIhanf3dqrYZGA0bpK0omvVYi0A
mfKelZymqWC2PCHaStEns4vg11IqGJWqEHv4dlaTBovA0RzVwzpN6BO3uBb87C9EwgZKd06tEcjw
9GpQDEhkE2DmjrGt15Wwq9UlOyDGJ7geHyBIFmveGTKOi3D7aL1Fr1dhPRf5xjiM6jt96NlxK1Ur
/IJ4GUdF2tALenwhG2g3Dj0zUlZpqL22LEgZFjF81zRXkkaEnPirio0YKX5O+aqfWdEl6e1MX1Ur
vRyJKpc+d7YryQPBusgckvYe8cuFKfTl6O+uIse73l/8JYQQAP30SXbXi/BUC+8iT1LeEolqwINL
JAp8e8tjyAA9R110xhgC/kQkdGVyo/BAW7Zu1ZDtXW6PgWcT5o6oWqnOzNTeds41uAKcHez+pg0f
2jtlf7y6Y2+mObRU+oBDdU+utVhz3uPPdfLAKYudJLKZZP+GGOhxHQfddbUCWkYTtAjRv4FDXPei
IRj7cdmUWLhcYokhnNQfzm33raeZVvNHea3Ss0IeMjt8tcnCgVxp3mKqpd2hhuAzcDslWaJ7fdVw
tt5FQtsKdBpxIY7h0lNlnJqR6YNQmnCxP+tINsZbG5D2Pd5NE8Qh/b1OBEqFxhJe68V5/8UtFuk/
piMji3HJ04I0RC3en/vW+VebJ+0ihxCQq+TVQfNdIHZyxOSu9qRejSIyb7Vf6flwesHp8z7sMA4W
DVP0WZ+riRbf9+FFQY4lY4GnhAVgFbM0HJr3HSCM7EvGovPfsn0qvSl16M+Vkb1/DdZgaOiIB6F3
zXZZiq4lMj0coWDvxkJMQEf0Z2W5rd8BytqisJX/e5kmbH4V1jKMM3p4EbGx47/2E2Jyh+8bPbIN
tSu3AYtwUtAlHNpmEwDUpMzVXxuw88kgalTaNodKG6bpX6Xm6dvPjYcKsfokCkKXqc99UrjbZWaw
ZfOFyJ8lKE1IgEp/+2S2FrKqViOkX4jYB+8SMCLP0Q3qCA5HULK19ZS53KKAW+0x33JMWT1qDXss
DJYhc9u2fj4xDoUnBAChKTuXCxqiUAZS4Bg/kF3y8vLOxd8SRULURL/hILE7IgOGMlZS33gdxoU3
+Bog0SEhMvrdJWxRuPUsMoz5IxRQMC3cI/RjdhLpYNDkx6BDZ93GNPFHQzJzhp4SBY3B9ftUXydu
VB2dxisNOxG+6l1gM2py5Ik386kcacJW4MWMKLvMx04ZUb0Wqn8FMsxnEmWk1vsZMJYn7r7tGWG/
bQtkDPthuGcK+dOAhbP6bjmyXin/crXapK1ZMIF5crAgx3MXIXz5ekz+QSSwSsvhbOxKUgAvwrVu
8y5hZT8xrrdjb2wvFzErgGZqMCpQD1bvHWgKCMpSNVdp+vObq6xpAbrokEje9o5MwCjI3ji/bVz/
LDEjnEL7I79WIn5t+CRgmnzA9Xh0XkTYIDGIS9wsBVc82tAxOLmsGrkNqKq1yXRZXqV1CbaHbyi2
b1MAdMD92UfgO2CWVPdk61O9ZDN6+HrlgU55TjhOVCVBLq8oAYmC5lGBIKAqLlJJ12i+Wcjh781T
rO7c7ajpQedm1GRjnMIJZ4GYnKC4IR1yrx1UpWLuqshlDT2vQ322CqSlqPvPKn0QYMEKuQ4htjsw
s9cvDJdX9kimMmMoQ5fZqPPS6psvR75hHExEQQ6gTeRCZxQZonqIVqOKvYIKES+4cI/si9LKIH8Q
hcnyH0WX0kdOr5pw9neTzu+nfz09lt/ukc8BrNDExoQVtzsww5u4MLPI/uLl0vtCbScSe7O4BiYN
vTrthh2fd7Ukai+r314XtapuoWDpRs0db0hb3VOq2Q811bPAsf669yzkty29zbZDeY3se7rQn16J
469oYN7efPd8TnKfzhxtreL4jiMTy0bFntv2dwGVRzxlsMHEQrEx1HNfplnJefmDrhXawTBI4Fru
Mmj+QGqI0LRnz26He6z4lwF6LClZcPsWPZimonaaSVusat1axZLFhyXJNa3UnmvNhxeQsazmLJso
yIA8FTuemP67NWhxBHM2JkCS0IOx/T6Uys16i4gakFpV4Jsi70SInl3VbRmlLQR2jTf+IBPbmGrp
yX+TbUzdZ8L3IDDn5Mc1Td0lTrkZRrjjBF6VduBvvL5sckAdV9l8OxWvkD9T82rhI5s/t1aiIzf+
gVAB/TkyNqEwBoiAYA/ZoiuWPlP/UKQik54WXmfacxfuwOEU+CAjSfs/SEP5A10JZnSWS6MjcjKd
YI4OZpDz0vk/xcBHg0EVoIrXAjd2YZG9GKhDwzU91ZQPSqO6kdDj12kk6XQt+B+9w+1vH5nJ4eNr
KjBEmFTdLXpbsdkDX3speQMvXAn/3CJDW9FkG8pXPIBKgsLBg6Mxk62Aa85SHcY8z8RnOz0oKHY7
J34eRWIEoKjv7XNMR/SuapMPoUHiRKU9XoRbCZi25tSS47PLNYVWi3BylvhfOPzH5ziF6gyPYPHq
vH/pSiJWtpbMrf5Lnv//tqyUpG/fdOps5KN5bnDZekJA7C8p5zZ/9/eeOpSrOyw/+jjl+LmFnyyE
hBzchM5YZIzicaH1kvzRsEPqu4G9FuDTTNMMMdAE0ZW64FJK4sCqbA7ov0zCcjQvB1ZSN6bMvMMo
cfdfFld42niqS2bbmE97kwxwPC4dfZgym6dqFDPUh9wglDYvYqzUUYM0NaQYKFPp8ZDtOj3WMHZv
8D9e5poznhmGQwfetE3loRCVR25Z3EV46CA/itVCNik8Xx2hjTHgn8q5+5gMTl2qzlxiY/T4enAc
T/oJ0gZfo3xmqKX+7RHiSsIkLqMPVnAr+kHLXphMU8MtjrJAuG9qNBvLSr5foR6eZ+mhxJb/y+Yj
qpzGNm3LciducB65rJUUmIQ0epbvBrB81mDxtbSPM5Dtxnv+vMLaK1L0uUYrrzf+oahCyjUWLuwA
7f/Skpy74o296x3wtVzeV2mjbfjkjAfWzwmwfmKdgs0kc63jhcYAQnTbLczziji3JYgvIx55KfrM
Mvj9mlsnzciURrtlmGiRerM70IKXipd3EmbSPUOE9fUGhr+iivOFVUs5gIH0joddXhTFPs+6u6Lu
6D7x9eSkrnWDhkN8Y5cNS4exHX+lmnTJEOefT+LIlG8xEj9H8ubji1xhMHcJr7lqUB00lqkGz6Lt
w8xyAWE26oHZWR+LHkoTX2tE+8P2XfNpwPnFjYUGlX/z9cjoao3L9/YQ2GalG9oB44GkHlpfPoEx
DYZ0g7OTb6hi05uq9j8sPrBLBlrFD6NQOTNUSIbRy4i/5cM3XVFN7xwqwhxWttS6+wvd1Nz2/E+7
aQxwkxMiLOj/N2DoeIuC1TQca+WPHKXDtz8HLio+gp82haoVSbzaKr2AXLi6gdI9YxMT0MBBkvJI
5Ba5Z4+hDpUCj2AZZY1nhm7GsJoaycb8lLV3+a2lfK5eRKqhJH0HB7FLv4BdKes8y3jleE4SqkDU
AwRHLD1P6exunw7thiL829y2+yi9wuAAWv+6vEE1ZgC2LoSK6KXmhl1VstkIZdk477QfzbmA5823
FqJkXcYzxAE/OLLPHLqgtIiEa/jfE6n/owGHBLmRDaovQYybKi17XEHum80FE9OUfYwLwwvCVqzi
UI81HgAAp6ZwPkbshOhHZi83V94hGPprKi3MDkGZP+fYAiuTwgd3B/jsNGuAS7/JnSX9OIZ+GaFE
HPN9qyKAXO4+wqgrSaz7F8C7LskoTIaxnsTrVWcACcIwhI82fvGh7D6sRUU9fkdKghfd0auICNDd
hsbieODrHSizuUGdvQNH4aNlM4Z9yl8eyZ2ZrcD4wB+1x7Qt7PHE2ZC3UkWCUDDg/49rHYt7YI8C
NEqKtgs9s5TOW0gy1gr1FvAQE7e6DybE7LjfCnAdLAGkxk9Q4+Z5gNTjr/34+JnG3Yf7b0mZAKY2
ChFdDDj0xD+ZUac9uhNpPmQ0eov+hXyWT614BjYudVImdFBhCJjPfBx68F03bgxrgikW1Z2N75LC
TsCNE8L6Jo4OH3ebNab5N/skr1zxWGO1qfRK2lH9hrAspqwuqE7MS8LSAQ7XrvflbMFRBCVrPdKc
8u5/69VOGY1lvyeFbiDRqEpCY3yRkjpQMKr4Xtwz727aQFhHyJcf0P/WI+/EMLZQlEBL7XJr00Ka
mmBrrP2k8jf8RsZ++eD4drHuBSwiEjyD2Z/puXkRXuDs3AGS2Nvmkwh8ljCdpbBWRxDAzXp3wMXG
6hpszQEXty2j4f8JRvAyGUSrV6r1yNTzq4Em0DJTM8rDl6mQko3mjpWDYYMwrJ0JNpT+iJE+AJt5
6lbpJ3ZgVYKVMQQhyV5V9wXVe2DAmqacgFMQ0nEUkNLJhHW9xBWxNVajQAka8yEulDP2ckNJFFji
LNJUugmXt3p7MOAtbRXYR2gYBhLQD4O+kIhSH1K20vT4jotuMN+2lmqrsd+TLw28FaoHHE6mTTfD
5Na/fcnstQlRzL610fM0fp+EYYSy2Em7KlxOh+XwGIrRzuFCfM8gFMwssMzXqqoty1DtrpNVoYSk
uY1NFs3B6dwJuUt0v5UT/zavd+oMBmyONPtLqSM1RT8Vwhdedti/XgZcmhYpDgRJqp2RkkcdFIuB
veU2XhtBOEuh7jHN/mZtSEqtN0ERqgLozUVzHrlE4sHLbOhS8jBRF0pjciyhgaGN8IPM0ax1sCEl
QdQyD+VwIsqnPoAGPyIepGgvGVaIif0bfY1ez/bf+SlGqqyKSC9eTQKW3oXI2hv1UKUGY+rdxT55
PTfphcRojCqb+U5w7fnoqu3yELwbBZFIy0PhlJVfEDqonaX2bd3oedoZTcWPoRw+sdTH7zANf2ht
OXj9219ypY1znu5aH7M0a1LdR8VLYS9do+3B6/l7NW2u7dbdKb5Vzxi3d2cyNhUU20a3kE8KGLY1
zzY/afUhsWbW2/Ehgg+toikCt+TsA/H/VNgC5WpsAn251Lcb/tOuRfP0enu56jdj65hM3XuRZk6M
DnyndFMrL+4xuyiKYCojShELXsilMDjqANucxrOXo+xQGG2rcd/Ksv16K+k8/Gvlc4EvQG/63mbu
JHwa04lPrrqGnwueqxhUy8c1XMI3+Vefm1hPxZdYyNI/AivBjzsoMzJapV9Rw/V9pcJr2HqhpTDT
NyQB0Qu6fBC+JEd+q2MdfYwUbHGF/s5eGQRA9QlAvrM12g5irJRvATkhpiPyZ2bTEliyrL5CCdzw
YaKoXBsB4vWpwgJaJnB0xJ/fXMN6YMTlLhmbb5wFKdBjdOpEtlcYseXOd7n1eu2fh48oLQ+CjZgf
0KUSCNrXu79KMeTjYyA2Q4BOgb/to3LASyukieV5+BlNo2P6uLKjWyyRGbcIun5U8lDqJYwmiJUm
+tnUbs/vgXuf+tLUMsGrgVLVK603aE58ixEAljZex/oAb4lMI+EPRFWBzTrBJLPYQoT0fOaMcaxV
dP+MNj4NKCooXO112qe9U7Ulz/k2obgRuFfeOwnat+eLs7Taco5Kpe5FskkdQDmaPeW3cj8wIleX
bqriTTkh9bZ/667fUdIyynl9rH8keu+B5r63HEZqJy5eq+3Tz9icbo4RQ0O27Y57q5AcRwuOHLQT
+kssaZ+OaodOxINblNnlYm8FRZiyK1QX9xM0SeNV7dSCUWybca4PH8eZI7oZi/2xv/3tjPOuP5qk
W6iPuKGX6sAyd3jmRfjbG64n/ZOqc6mFGakVQKkojGZuGdh2AttlQmNcQH0hpuhSjJJiCX6NeIbA
HBZ5GASfPu23h0pOxjWzJOliQ3FHtfOcDJr0cRDxqizVmArTLmS4h5OcXAW/RNO7LN9mFwRWcpLC
ZoM+PdIVsv7T2C96ziHvlR13YPVUAofD0WjjiGyntO+cNaf0wxX5CuFmWCmRW+vGQXPIx3PfeeMM
ng1GsLMKSkH/MMkXZJQ36ut4lzxwPi1C9tze0ZMlIeDskyP/i9n0MADLSRk/9SATSXS/wUH+vJtI
Jubq05Cz7jl2PRibkyGSyWbr7LM+U8eSYamvlJyaTurTn2ctC5Bda5UGHqnbC4FPBEkIS+QRzjX5
yCxBi8rmkvLfMVTlIvOguJIkPrhlfFW29q9BJpcWJFGRaBhk0gtPTW4CXr7IdPTwdM/XtQM2JHg6
h0zqRsQ7KTnyz0r1PDI6b1aFz1rag1xH8DsEuba7EEUjSFP9KRMUnAEwZUn7xrWMhj4Aq8RdO0Hg
bT0Nn/AclBIMRqsr8xtY1RzrQ1Y9xLr7tq810YcIHgy5NPLbkNJj3m9j2k4XhDD/Lc3e4xtrcoKw
tDrBu0zZlyUpFn/Q47D4dZAz8g5GP34/15rNezsPJCIi4B5Akg9B7G9FF08P83jGR5fSSj36Umx4
F9ZM07JBDPIzLPqrW/hSADqhx/21U5D4pyAh49Pr4aTLrc0MRlJnsYLytYGo7r7kN9AtHuDnU01i
LoDtCs1itfu6YawsmxWxkgyc3jlemqJou1tMlBrExRphU7W6T8nBKRyJCUHimBD0rtbajXoUwxqH
tLyatYVAWLWlieSxTRDssOOg2Iv50NwugNqZh+eau4tz7aQpwExwAiCdRYwHgBuV4mZM/eh83TIz
dnbocRjvTAx972NzH1p9+bdSa3VkW3G9Oqd8uvp8NS6BOJ3Rg6SmqLovPoLA1cbJOKYiRom+0hkb
NSupfC4OszfYC6iq9l+kZQLhgCVM6Uav6vlSX3O7quiptzKOm5uNAk8+/CoNHv1ATgDyZtMQtyPt
pPYGcg8fa5X/SO05a7QVpVxRFvm5u7aREtGGmJzg8yyCpENFtzObCfUaRxyjWWPa9q+MKaAN8uKZ
VK2lqVXygnOg5JTAGi8JcrlpkwM2G+74ErFk4cfwqGJUiDX3Yr+P39jLLECPF1bdxr4R/gOL7jnP
ogmv3F1HDuRRvNY97ixPKtUNfPjz6nNuWDTS7AboHIkyj26CR1w6FHpVObH5eh8ymbylspKgd8F+
nJCp0h2l+cgeiATp511m9ROpe2nIYT0sqlaYCqb+2JZssX8eOAGCp4Wk6Ab0xTafABPTj4DXCDnJ
b0TaHX8jbsdPF63+chCWW3X5jzrVLEb6rPAWsN/XgUS0BrXiguL9ENccCv11+YMTPH6lSjISXy0h
bgWIq0FuFBE2HDs2+yFgr7EUrJ4/ffcWk7BOGcRUp10V8//0Cdtp5wlzYsTBx3DQVDxVskrp2TyA
qrRR4cyP1MJhVG6arTgl2SorBZIncBQg69pjqqP1OlKYbYCFQaN2Aptniv3EJ3Ei4tnpn7xs7DzV
QzbgXT85ZJ7mWBYHksN8SFcr8JXZMxFKdp82IdTvF8uyl0HuouF5DI5TWGG8DszlReyCDOzV4Oqe
D+13JtVv5bbH5z1sGryOIFNbILq1R+3kUQ9SshQya7y5fc5BtRyJZjL4Quu2R13za5GNs/A/EWJJ
9Lh+6mjIAT4JTWey1AgL+p76MblxcumLNOFCQmQIFDvTJfElvxgpP+/cyk5MRrEVPZ6Uvb6wJQJh
mHGZj0axlR00Q4s5hTVSOeNA2wYkWucWQieT23mEzl/8gyw3MCSlh6PwBYxaJoMlg+jZC6Hir0Ki
ZA2fZKwXEdMRqiBccqzdiFwSrD9vIsnjJEXDs82hMeBVOsEQ3MYkT3KYBfMauqw2uw/gGKhd7tPg
WFb2Nr5EHoD94v4WOVf0rHIkVfmVwkvdgydhnnfhO5p5OeFHDFJj2r3nh5sgENjZoZJtINN9lXV3
nuulv3m2sIc+f3YFCAeQI4NgZOg6m9gIoNM3QDUlcQe0KsQqrKQwF0GIxe0s0tu8dXm4v6rX+GcZ
L717of6/pXb8uA9PzfgWTs5H9c6W95Mnqm2LVig8GtwURc57hQCat65sYbW4DwXyJcfqY/9jQ92n
OX/3soOa5X5gxw/Rri7dt4n8kqm9nR3KFw66xl9P49pfzJmvST/1NHeYG0pDNjHtUCg2Q3CBLyo1
h4ocA4wMS5Jqerm3Esem7OfR55X9TAPkERMufCOHDJgsjN0yR5gsLte4xfJeLTKybez12fq1wyEy
F1PSnfiCfM8u0xxH/FJJRb3TR5Dkq2ssDwCx4Zx7ozwcq8Y5lm6yPJHQ2SKsMqBdkNwXxp+X6TMP
fVwx1rY6AyTRgxkHKZfaolhqt9O8S6F4JnMEV92vmbvqZQ4I6Mi+rwWHNdbH18wwcbkvT9Qnfhwa
GqTWrnuMHyCNPpoChVCha9YvY6X34IE9AIucmamts4jvZsBt8kR4yPqO3qTsa4FJqaUZjfSfXrrS
lMbuNbAE0ql4U7cUOiGRjbYBbVw52R7lMgaWyc2s7K9jVuP24NP1NjUEw+/y0TmPyNjeQvRhjhYt
Taf9FUjIqzOVs3bw1t7wXF35+4p9EiNk9vdc70xlo3HXt/pNj/RH5b4rIpyMhlwox1EXSnPOnj99
0JtWpeKG7yFrxNhe33Ykz4Lbr7LfBLInPafhjnbAg1GZ4KZgOvCV4ZKU8V6hiWEuQRo+oUiIkrBr
G2Ag9nRCE27ab6mhfwxPhz2njdN1Y7Dpif2qEqBCr6RYlqHJWhRQmTfgUz4NPXogS1rqRcIJaD7c
brWG/KNUfXSRY2VBspAnI/8ceUcQZ1vplkoBvElNCv8XDEtV7s1wrWE6OBS1eRfCKauWiCwD/Bq5
1Rsxn7Y6xXDnt012Id0bo07Tak6yvUAgbezZsZy4SvkEA9C2QGpABuudFb6VHR9tZesAM8UPIbxH
Y+4evJe3/ABSqh3I3ulr7Hohcetsx1EmwWgBsEdpXsgWOUqxSuoYhkM6rCSuJ3BGvB10wpCm3nNr
wKvsubZfvI5GAeJ0m074Tjx5UrjmhrUrDQOGDu6Id85v+ZDK24JaoA9OADgRjuio+RRX29HeUchR
23xgrp++a9tQQ2rzecCfIXESeebExfHncJ3RH7qx9NPVmZ6WbbmVcsinw4GMe+FARDsCwSbXQ752
E5tLaisc7bnwtTIj6BIP19sifXyjZZtDa3lngLLvQvZ9LWNO9SyHzLD+CyjU2vQZKJsouKqHulxz
OqD67iw9ST1j6V8AIjHt+8F3gDCOhpkR4qpC8PFowFNQozyVBgT5fCj3k1o/hg1HrbQUmtPHFGtC
l/4lIgyuuLVQxp7B+mixmA0jSPr0CvDwPtTT+FPmV+GnvHxajJZmzi9ynU0w0Qi/uKygvEvsebRV
8Uct13/FsyuqmqPxfS9AyORziOxMKXCxrGKhi5SMF/A+7ws8QZV8n6f6X3A2bxZsm8vFeIq2iMoH
+kFFxalkWqClNntEX/wI1y0Bg4OnOcEom0Iu0iSiu1SlDmexYHEiPYwoijNZJaOgnHuHPdpqybhw
tuO4X2eGwsnYCmtYrvRrNdMvLovwtOVQ/PpPq7/T00+6FtXCbEhn7j0Ib4d3c2ov9fmkOYzyQ5+c
TLwqRiIgVTGZPRs+AcTdrk91ICfmXIOH2LoQ3cckehZ9eetizefOB1i9p/f5Yi0XVff4lHN0si2t
e3fdPNSvWbrCJwyQ+hRU2keyoxd9vPik9Q+J80IdV3n02ZwzdqlkHdo1v1t5JnPJgTJG/nmzknN8
z7bfJaaj1By6ees5zKuQ1iBBt4i0x3xAqOyDnFP3KrNYNp2nZ/aA7tg2pfpxT1XOypLhrt70E8xA
9yQ62/jZOumDzMiMKbe9LaQ+A1YXYcAv4KrqRmvxdlEfQcyShZ34f8/iFz3NmlAxU5IcMzeE18np
JB+JOGyyHRiw//pfwhY3IyBWrIjl2otXNO2WJyRt2gJszwCldLyTtwptsv/wUt3sNaxHRsEekqKD
MEP5cFUYUZcri5hBNRitB/WZq1UN2OdzBeKmICIqFjlbTc6qb5h0BlGjWS4voqf7+0Dk5KuX948Z
LFNwiCzScjsDc+xgqEl2arXN9+y7WUClnVK+YP+iUQF0SGAz7F7oR6xzr4fgX4fNMpB+sF+xn462
UVwwxj+LQu/XE0ZAJxc3nnH17X3jEfGKg8/IGw72GMP2ji4KqDHWfyrUbgYw0eOfPrVwWBntuS4O
lnYKtsiyZ7dBYRFVyvm6/ypMuY8wddTomR8SIqtKjB0V1UH95pJVXtYdYq1lhlqglahFtYPNk5OT
wTTkK0DbV+7mSWyoOaaIGZGFOT6AUIl2HpUB0RhFw+8QGnpkAQT60ErpAOjVbW1LcAVrre/BWeaK
yVeDncrhASKIfgnAQHJckUeK31GOGL93sT+IWBnpZjwli0rVPg0oYpD2S8Go6B/OgZgHiknBXWVP
9mZ2LVoAS/TZUTpwcGpMFJFZIJAAtEmyyAtD7Gs5pE48JP0n3tW4s6HEYiYwIcXPRpL/QLa2S/5c
kVMJglV9OZ6m3wk3vujXz4+1YNH0qGhj9taKGAVAbnTXwedb4GAtHAf5rJ+6EHVJ3xzEPnbkfXYh
1HeYtIPZ2RueBFve6sh7SXeLyOTmZpS8w8GgqXVXUE46HgvSK539ic4kteXPMNaLrRcySV/du97R
IF48rKUypXvkTJWQe4UuUGYGRiAXHeMQ9Dsfjcc0KFAcrY4rpx0gmmKuQJlKxHwvlyCz30BW+/RW
+/R5jh+dByyJk/6VosEErp+P8QBBqHoIsHtKYPUAMb/f7YtZPSFK8leimPpSom6lqn2MsLaxRTAU
kGH7QbGBxHBO9ED0NY9zAzY8M6HqA6M7DTeaVBwJU8mAZNG2P7PWp7sRpnWtYSuU16XYpIsFE92/
gHpgd3cVt6j7UDFRtcA9R7ZnKS7XunQvdbIp1vQH1IdofZaON4kY9uMlBBp4vkMZ0uM8i3isNKha
fhiLBlL/vT/qsdL9Z3b5TpViwdFcmsik1IiEFN9brTiwt8C3CJD1WfXfOMdO3WEOuuOCkDwj9iaL
ybCDN4uY17H75ZX98KNvID1fZD6l0Jl5u+ygaa7PbELSrQVAFHcy7lKMujehMG5rvtpTa7wmWR3J
mxKj9LNeBiK1ZN3wDq7NFejwDxZI3CzlOn+SfjxJsnXBLFcr7umpKbnnjxxwnejkWoK4pW+TJ7Ql
G7rks1MYzQnD4QMx+dNPpWGOqLeLxL2m+rkKcpTNYhTS8r1O7CaM/qZCdpvnl2MwE+YzaUQjc9Zi
haEc3TIrZMfSqQ2rNR6YM86c1TNq0r3vmDjLemXJ66+Ote/pKGDbKQ9pYMRTosa7bFbbrBBzSfOx
jWRSsGfr1IN+jwoPfA+dYBC2xUSsjC7nNg/feIWs1CDuxor0WJOgmJLKA7DIqIi3ZOdWnaZpQI1B
jo25f/LyP/1XLOqQIHNI+gzMDcKJr6rwJEQ4x6f5dq9f30NGfAgni4Rq5BwXWLN7repyVLsnWwnl
6gGdRuz3mSxi7g1x+Txrpn78nxfEIKrR1kXawZj4HecA4yR+evWEfHizdTRk3dnbsoJsPizvVoj0
2JR543dxfY2nwFF4g1JtIAYXucNeaaviVwLQ1dyCJEDNrLccB6HYWA3oGik9zcfxDsIzK9JkIyl3
MMdL0e+c36rm+YRkyQL92HynPT4iAgzd+NhVO6Gc1efUcfEfzDTodMF9gaemjoPUDn7RtrgseZrP
5b2lBBSqOum0YncwpqzKvaykuLbfwZqtdM0EAAi0zOkat+envMVkGSy2a+3vNTibQ1ysIvdmXdBi
IoYwB2M2GYFIuBw3j/qyBMKn3xs/A1vkIhwLEe70aMHWYIIKH7W3dHpgHKDaSI58qh96jBGrW9Uk
HCotSRSazINPOySV4JBDMru97GcxqmUhwrXG/zpLs3GpSGeQDEne2mbP3X8e5JRjANNKXL+/wjQQ
eGVnlej8214e1Gen3em9LsvmxUVE88rnlYLlOY4aH/zQswkbA0CxOnMFwuNDhFDAkr7A19I1YI7h
v+uz9IvxF0Yyqupn+vo1lyNZXfTU2ghtztORxTUEq542MyALb2a+JXqgiw9f8ZYJbtOc4Zm6e3rG
N4b1UZulmeWFM8nGNI2acfGN5MjXYvjtly3TUjnYsjuK0LmZ/P6NFCGOkx8AGCpdKw5ank33cwgj
w7+xIkOx0ETMg1lkH3/hQC6skUJIgxZ8qKeElV0javvJBHGMlyQy3HXul/X7DMSMyTuAdxU7Iqh5
rFjv3jt2RiHAj+yhpXMk+BywmruMBSJlrDtGBT8nvdn/pf3Dp640LcCDh4eGkFpqOJ/pFK0gl8Bm
w6q7ZuXbo7sWMUxgdAKphOF7GtvknjZMNee6alhH8DnaSElLw9wj1wb50rPi/gXl20Y3USufUs9a
bO5wwQHm3AslO8ysLzzjwWMMEgacZbAnL0kc7MvZrNtrmsBV4kQVfJOaaBqJFm5UkI4+Sr5QwaZN
N8a74psl25iSkazCfTic/6yLqLT658yJKc7agxMfVtLCWrhFh63VYodsRga+SVv6aRLGxlYIVhFl
4iaSW5Zr7dqPTgth6gRyy47CfLniKeAy3lbIGSHyqB3Q8hFiyNAoh6LldzK8jCiSSjAMN+xbkfC9
EHDbfAWIJnxIhcWxmNfTZwMl0kQV9mMGpmtav0rtMovSSWGG6YhieQ8vDHdzl/ZO4Mro8wn37YKd
x+7p8dSawgSRwyYWNk0SiVOluxzI+HtgcZt4bKPJAIf2n7RSvBhYhlUA35xWUrr9NoPT48rOrCx8
VOal9vTl9teaO6Xr2jv7mSlLduJVduVKq2CtWy7onrj26mGdlhXX0CkNtattN3Tp9rBBYm0NmfU3
RPG/hJGrFsjtDRTRh/gGYCX/PkYLrMCfweFg+zqm9et1uSoRwhSo+GtzWWHrtcUZ3b9Xkt1FuX2F
BH6c5bbBZIPlQQlmNO7JEZZQFATs3RznM5IPFZ4dJsBX4ZzEgrcJ4gyZmvalz2THj3P5oDItOaIp
sijj/GZwl5fyZ5/w8MVrgchcxl4MN9rYbOenSakSSHh+cTm/G99X0cnAfJs8otc18ww1YNmJGytJ
gOjeeHO/C/dF9kgW5PVzBH8whzfQLkQVSweRtI5g8mD+98zsPGm8M0GQOrllOl8jY8l3lOCTKvz6
S7cQSkkzjkDgAX4au9G4jm00X+kTLbRYyc06f/R+e0n0Q4H1gwHnmPd7xP85OfEyoNUZaOM5DXfl
c0/fGTnxJuFiV5c6ysG1jxbwq/9vDULq+aDHoX/kxWyjvbaGZJKv6PyWspW9vn4kfEpKR49niT2s
vGk9fDwlYrWWec5ix2SY6HBR2z9xPU5SFwDhCcKClkfhmc5+cgiJmh+YnEIXGCkAt+YFjCsQZbGU
1wdkaL5RS2DMvFXIQUCuDWMeZBiJrpltJ5LfO1SCFN16vNr1DH5uYOci35i9t0D08x/0o5llg+gk
eguEgc84BkuTYcLY5mlSL9qwoweTpBcXTMkP/oDTjLLNdkNOX/FDqOYVcnMMtAXEoFFEMQ2Iqr/O
c7JNkYL4CWsuflcuN+lKpkn50/U6uC2ZVZWA5Al4Zu3gI8J/2e7MMaYIDAYxkOO2iOPdE7zNr2uw
CPn7KxoXbMBB+Q5TuMBf1iIdIBmadZTE6IaRQdq+Yzg8rj7sWDg0DKSZhFXF3hKe5e3MBaFbNkc8
WK3ESI4AzoOBcBRHN4WlsHTviMZXdYbu8tJvUwTIRrRy18ItGdi6RgmHnM+cO1uocgT2b0OBVgWz
M61mgTa8ffby8XbabmFB/UZVSSGwTGHgDRUHvkK7Hom+yvCvqscqq9SazfbqbEKvdreU9CvhwvR1
WTBAicQ8TTQZqNr4eE5Sw890Z3cxu2F59uIOYXGRLmY7zC1nrtUjlQ0nSn5pHu+aUimfuaD8/YST
fzPmPaWSqCnqodA511YBzvtP3hU7hj7SkuLr6enmjFmA+WwGwAnz4bLiXtKEGItTPRs4YT4cc6pp
8NcQbPuzI2Yt7ABIemJlizOKMz7x4Dg10tpaVb2+6XOSYfehTGF0ALPYTlYtucpUWbom4MxgUmks
eAg4fsBtxL76aqfNaTJwtFhEgd28iGG7JtsyKpjhklm6BqC44Z4CbRnkSEQzeFjhWNcCsriyr9oV
+nVD1Wga7abLOkoV3I2QDT5mWiAkB1wQfV2IhbOi2EChYijGgLESAIcniqenHFX8ZmmyP+/Q9SYu
Px8aGQWi+AO289Aqth5Xsu9ZxzFhPlYoGNtdxovA3p3s4CKbBEXatW7Ak7qW3xNQ2eX5haQ0dOwi
vlfzxveTFSkFFtFrv5Md7HPcZBMsP8YzAJWXhImKI4RzDIjEFRU392idGheOei/uB847u6/XFP4R
54uHVn7d+fSdo5VtDjUFY0P8KvUYACP3hulrSDkGgFdx61/kS3FQyR6RDLtxvo4NknVmYsIbCTYV
JMJv2g9eH9Ew5IuugxdWSSaV9GehpNI3Onjp9M6dYS33S8T0U1HylC0uULZa8TO3r1T9dRLKEDsa
cXkxpPdxNV4MqFj4+VQBd4xY5gfZtLxYsIeoxMPo5Nu1nBJi8rF+85TrINqEmiiSrW7cmdU0NVCD
+WdFozBMgD/7S2IOyB2+dqdtdloUDPMug2FuFFmqlfXue3Sr6dUApDWM+RwXdoEYKQ1wK5ez94Tl
gJL2s3jZnETlIE26AGm/TyrVtRl+D4FceyJswmCa3FNcXuBsjZS2wya4ROE39ldlBySdIFK8218d
vhDUOm6W/FaJDs/+o4vVf40kCHfDFXgsvVVpbUXRI5G+UwzOxeZKiauOcXo/qoVXz2g38BXWu77+
FE00iX/U+Ny8ONc+bh6wzpT/5QK64zRXbw4yk90I6bogjTt0bNqDs1/2uRGmTcJl+VXvfoZQaJEh
Tbr7ozIOHFl+y9NepLr/dwyUipB+DcVrKU6fADiWi0pYEGSlV5md99veDjyxAxmaMsQ6SayNkbFW
aggFszGgHooSnI051tzuDMLjU6ObH06Jv2s0cVi1OWhDviD8FtRL3sy2ae5fr0WGbqyZHXvJ+XOc
edlol7RhOqgA019ctH+qmTru+RbzYXaQovIWwPahHuNIhkMATw0MdT0Hi55ulk3mHXM2WS4Iz43r
XoBrbLGR+PqpEayCR9k9PtcHyOPIJBRE3tLUYQuP7bmVrhUffd2JcZ3zfMwkj+BXislvXFJbFtwu
q7N1Vv0mJf28jHvitju0ZyBqZmRL+G8HciY4HXzJQNbKl8y6MvfYInqJuPS4b6BE2LTeILVUuCal
pktTybTxgINVTpmhw0yzsR17J0Ut7FP40TlEHuPTXx/xRb/8398o/zpHAmlqyF8v53xcjMLsqDRz
UQwCl/715QBm8p0L2ksmmyZNTlFTIqzAeJ2TtdwS9raGna5+m/bf/ZCgLab5KViL03Pj9W3FkLpG
X1XkmGx0ilFu7lPh94gxoirS/Lfp5WDVnWh3CcEsrQ8pJLBPmbfxz3J0IRxCnMb2BMr4fp6qR9/e
JY/MQJaGXPBZd8N8mB6mUNAFqMt01DVw8Oyp01JFubCfUM6seaCLwE3QIybnDaDNwX2hR1Qku38r
cDemULg6nBktLSXCEYPb37QucY2ti0T/6qDOYED+O91I74O5rLmQQMSZOq8D1N0mlRcCzHTmBJzV
1RUaErmovAFvv3GKnBaD+qfi0z3SvSG7s2QaIE1XrCqM6Z2DSMCQ/bSnH6j7RTosxEC7Omh+hTkd
EfYwiDuu9S9h9LH73wLioPShlwIA706+RvziAvheRbcuy63Or4Qkc5LFfmhMKo6klGeyr8CWY5DV
Un1zYyRwDdNvnLCnxkVpSBfXfqsZwr+ET0eh72gPlUrz25o4I5RkH/iGOxKEKacnIlFe7xzT6QyN
VTa1tNrac3n2H/b3QoZ6iJTRPk9yuZPCuPIypyvkTpZwU430vkz4qmih9CQp8KkVmjmauTS1zKW+
1RKRdbDY/EvbBtbAc1IAkWCe93ZabezA+q0oKQuWJtZ6XrYZ9yFQWIJSVjitoazhjWcsreQGibda
p5IvWkIogvw8FPujFCLB8J35ZOUXIvy4xpiKogl83RUJ4LCx7ZDqrE97Djh2lbQwom/IZnivJAdf
sQi+rFYLbK1ngTq3VD3yt+jvRtYVgoLizukm8uRVOsbgPlBoAO7tCzA+ht+JxWvf7lkkzsONzM8k
2wFpY5yjdHywTkmumyD5IULg2BdjaBUXu+Xh63onyGoG6g+kZH7Cwavk/OZG179EDKG8RrrogMQ/
fd3j9odqQVQwVQKcbpMTA28So0OEmUzceOAhIpkHe5O+/Ji56r/31EH9nKiHZDRde+oKg2AkzyYT
ObJ1kLpqiPorslBeRkjxiuBlqW0/n34rOFtUSFq6ChRqqP8UTg4+tAgB9nLF3WQs6146bplTiRu6
lUAnCmmucZUE6PT80mngTYhUrKuXTqxqje5Gd4Jb+5wlm2lHWqj7WCnlwetwttWtKhCu+LuVSYiN
3h7s8exJtUKclqNDmpr5uTJ2YDE6irV8MvlPiLFndC9SRqT8AlEmcxJcRaqcFdugtMn+vdufwc1T
nFLCMrZ//rSIt9BejqfBXhJ2Ubf2IMoCbAmA2TQ0cbL/hgvahJSh7vDwDocoJqCLevLHQjdfaoSU
5TdeTXciyX8s33I56yF0sWpVMLF09wxHeDcQkaOVlqPU925xVI9exW69DRfwlO6Gg6nJtGmHANek
F1falGZz5uTolsF/eqEj0U9LPRuJuV19WyjwZKyIBSkuY4D0mLaBNGgjS1xqmzj94ne8GsIGdykp
VBALKYv4yxcWogm83s9oi0Y/IGaa5BWSpAwN9SCQ8hIVrdCtN1zrULVQVypDNr+YeUiEtl1ju5jA
ZYXcJJt2evLMjDVZbTo14O88X0tm4CTgJ3XPjrr4iz6g9LgM28Bu7vGcZCsfYcfKxgZU9AWMt1Rj
8ZcUwG3h9wQ0vmU7xoNrjBjD2UWFseoKtmZIrxuSR6aT/Ua7EsfDpd0btZSrRWe2h/qtjzlV9Thg
5VKGSnn8g90KpypD6val9AdBwmCGgdebLDt4jMqhBGyXhA1vZ+Cp0yGvGh4ArWV3sA2edDdYFeY2
+FAC+FhghcJgArBjMImpbntz5TEhHyQHTYbIfl3BSWaNmSY5v4tiYz+4lPHXf1kgvsIje76QblIm
FzGGqli0L7m9CJEGL4WokM9WsLTf+cEZ73bXEe/WVQX9fOdq4LKEW5e4nXzXDNaqo1LXabYjKBrP
o0I3dHERyENiVjtrkRQ2MX3LcfUcnDndCwh9/bLSuyp7zFwrTVm2O12X1m2MsdiPW1izSWTU4rBP
etM1YJYMrmQx1iZkDJb+xsLfauokC/Cj7I37t5sRTs6QbkBJpn3MRb/BiqI0Q67Ol0pLlNgy0/Ap
hR3iB4ryqxCqXM3I7XA4uT4KakQl912xWQatss9TUMcosXISMBEGSwbNQs09Nd0dDKYc3ZIsI0jn
hNd4AShc7oWYlo2q/tPD2bdcSRYXoxrJKL65d7GbG4jPhMIxJioRgY39+ttbgeLuLbdWzPIW0rKF
voKim7h38crs6xXKHYMYL24368numabLDHvApbqEL9YAWpi8CQMcm+DGCDP/HLey6H7zMMVtTwFB
p8KeDW6WCzY7rqETzCYonSbmp6MeEHiHuPNBzFjTYJuMhiF1x4t0SaJzoKzWvTwW2DkuORClTB3e
/3zRmzS0e3/AFFnH4pJaWWEWyKk3TXwWcvuwquQtkZhVLEo1e3sYvoXlMAhGxmOT4PIfXFod/M46
pshNoOGqk+Ivl22TjbdBCFRqC48FxM9x+iRlmlzPkLFJf89s4llmeZNk1BKVJ/FqIAm/HpRGOgfO
D1Wf8Xzoge3nMG/C0ykvNlF4pCzo+/rsiVfvZCGtiaLXHJx4zOobobolqGG70tnSMGBJUFUBG34Y
mtQY3B83EIeMhNs9d2dgg6q2ArOCPUQYgKEJ8d0dWsGZ05NmiICWf99RphcKCetLPBMMCG7RqslU
85+fc4CbEJpA82rXINA1MDzQHeL3eQaASJXsZEUAJTpzjbybUNHSoU7vqPXadZp/ukCyDI/V1tQh
V2xg6kWmHw4fUTrb3+F+5vFwZnUX2LO6QhfQqFCeX9NaZbSb86oJ5C76V+bsM5qTqf6Bh/cI4vsV
7Pp/mIV+Oib81Nmt+D+aiygaS2ill43CKqCEOz6BUHUHO1hofrtmc8Iwv0S4wHx6znNEE6YYjiNe
XYdSWCM/OZr3R8uvpFv2Qv/ZKr+pXbGklxYqVV0GK5NtOYWDWMzI6P2KMOiiJnsfhQkhGyOL2ub5
CwNxftRFR/kZbx33jbXQK+fWl+fokCqOEJG5DjbxT/WQW+rritcFsmf7U+xOVk5T7ZykYEGIlRaa
2eZsvAKPHP8SY/bvQb+yJs/7qUtUKTw8Pit56so7tdCtFTReiMdfSpdNYdG8mUR8sAZUGoW6rW2I
Zdvjx1z43smlH2thsb5YUNgnnsburDnyQobnFdKXSbK8KpruL5o36UclI6zbPa0OaM9nsVB7KUEo
mgpX6eRsJruY6kYWhmgcnNAX8bmnwsk9UF8PekQ1o48noLdaseYktk3UaTW676pn3fTf7hwCl0Tf
zKkXNoSNFSan75FLZY30P8opfFGToXtG29tb4I+8EDwccfAGBahm3l/zi8hDo2AT2+Vgd7MWpEY/
+ipfLLtAGmNsXXgHVwJwfM1BfVnZgA0XD+EV0/zQfKoEO7AXJvmrUCih18GQNG9Q6XGzVQ/cdU84
9qI71A+p2Dc2dvXwgf+hbOr+q+P0ELDMHxzm+jyp3AQJZjbtdT4pRhx7Kb/yN6Pu8IELj6+bhT58
DpssDit+Xpf+poY4d37173D/0CbbMKfbd6NRgk0ZjNaYrBEpR5HM4YuJczVf0xKYus4PAPwtHkFL
A4r/DWAGfP+swZwHyASXRQI4rCcm0HluODZodmKP2geugM/DjDx5HM3WKpb7Z+TIz6/PlQ7YNkSa
kBCj5aLrTeZNNpT3wqzqdtnSpeFdN7yCCHb/Mp4lcsDFbXTFGLKMRs8MF3ultbZw4z7YXp8HF7i5
pOfmj/MCaZQ2NcIPWEDYscdbaIBGQu66ZjnMvCblsY+gPVDf2dgdp6TMeCmosyV0gK1/1EL6GG98
5RUTt5380mQa7U/e5p3BhA3z7Dn1tnBDXVr5LjGwn6MEBcgkHqKM9h0Aej7D54QvoZ3CMJ4vJztZ
7dLPiq4i9xByc9orlagZEMKGi5Ldkv+xuBi14oeJfenFP+m2Ls5hP+t2XxExBZJDX5qmEZc8oQ45
DrKYeSaflIuCnhBCnekWrWCj8pPp3jKjVqvWpffEpq1Xdd1LdS/MNdlRJStvGMJXsKTPsBPz53Cv
088yDU9coqv0tY4G+qU8/XFe3VU3YJPKuKAhPY4+xLy2jjCjiXTdAhglkyuU4YP0kiUbAQ7mwcP1
ntCD/qqaYfKzYDMTrX75dvVh6UtBmELIWpBuYXkPRQpbC4VKjC00jtw38qvzYaLRYa8icYgsiBwr
v2mYqdj60IawfofYki0qUMOVd/ZjeADENYL9aAFpRjmemyG+H35gZj3L15Mx19gZxpF6wDR8yTlT
cf0CxMwLjQ+FulohwShT26xdI7oEK37GHdsU68DHHxE97U2YjQv+QkcNado23zW72vWOWE9HMWXL
nEuPXCY37+E/rJCS3+mmW4EYxV2kxlfAX4K54QtOfbFUuVYvAYuMYDVWbZZTtJ7hOcn0Q/luN4Zx
bfDYa5Nbr91gGdsduDV6gLaXOiSwv9Zg7q4Fyn93tl2xZzAbzddPM/NQNGIVWZA0pSOdi1Q+hEFM
D8lmh+fr+uq7oJEHtczslc4GzG4lPuaDcOXbXmXwlBimTesg5D+sxwWZXvch5X9NZzhZ/7HpOhlh
xxhMELBHwGWBxmKd5lBDsJZp56+DWyEO8/wE5B/GVk3wr7rTmf32x+ce8ZCMECiAJMd/wgR2bOXj
+AACoah1xpMi4IJMCZzUho82Jrb+RAhqEceZdrrbBo6OyqFVpDfJYtPG5M3u0kWevnTR6CPKKMil
dIb2tVCvIVMBpgzOWBrgryX+4UYD0RWjj8XH/X01773vuk8waq2XFwfwkwES5whQ0I5UdCX7UQpo
Ub+SSzgOiL+ReSIWdpoWObSC60uY8xJyHeAgMCeqOxlM9LklRn9bwiU85KCZmXoC21r1Ri03HCmV
nGPtqDr6k9dHMIWTP4DFxdade6cg0mipXAPxJkD4Iwarop4Ledg1RudYcmwzkuAKHCGm86IOFdLS
7SSoDHXlvJALDWlEmZbXwg9yD+9UlGnDrmWdvpk+2zGt8q4CytAgQSArOgI0U+b/523Skwi4+A9L
HZ/mo5USocV+DYl9maskq2nthlgFnmeD9aABWDwSEkjw0stAPSsekWw5/sOHuKXawWWRNLOLAbwt
kLCqVZfV0VKlJi7XEuAZvUNFsUA1jNiBVli+c8KrsxbP6J/5qebTBILeCBa/qUgQ1WRhmXGE8L8E
gm6nNn9WUqJV13kIGCYi6f89fK+lZ3sHCKeJDbU2StDYj08uYpTaRVBu5cF5/c7aAANEYBZucfNE
pUEHg9Bmb4Wss8FpiouMHrYqRi3r4YGKPMNJzs3vqXElYbQN3hi3phevWECbvLsk9QaG10OjKALo
NsXQVZ36zqW3rZLi0pg4fTOePl/KhYIOxCyDra2jSwyP5byYEVvauFJLqZn8Zkcih3mOj6WtyefX
ccr2+Fw5XrI6H7qP0Y8GX8wAyUR6tOC8K1+OUdgqvgdfS9JUdlnecxpQiMZ4D3p/uCozw7q/Cbi1
l1PSly4H6lbSeDSmbIL/g4vDupypYiC/OLo79rPB0fCXvjkDN5rj88MM5uHJMDnnS+UkxZImwDyQ
uCohc/Jn6Oz9+iN3ZfySt7QxBJknBXbccDFQg6JFWi0nhwl/edHwgtFtcRjSeCkB162HnADpPnMK
lkqKUN4/l8jakcXgAXrHjKxLNqkpgfh+3higkVVI9PP8ezf4VyzHXWl5toI5hU4CAVoU/QPdgxid
UXQ0wFjg+uKDefyZ4dWUJ29/jk1RQCXEtVf1WC3gzfRcr5puGzuSVF2Qzb2a2aIh3hCNfELIK3qf
aH65GGSgzFfFbrtx6MfT+AiQNl4YB4u2cD+QOUQVP3nSd6wILcRFmWJkOsQB1widL0kgpbfm8Sza
kuTYl1OjP6AWlW57uEY+6KkYvKnxxVxRD0JVn3y899BsbvzIfjU/E+fWj3+g6ws1vpqUn8A0ti3E
lvkZXjW8pbbE7GyiNacUX0wWqxGN78MuAtgFy7iRGRi6wiyZ4BRsk+2CZgK2wltf1mVWyj9tJ9yr
Ndgvn/Y4Hd6MnCDUdQPyQbBwdfLHWIj/qpoQHI0+uXRc0zfd/W1SVRpFDuI0+CDv0YV5YdNpa6Tb
/z0qZ0kzhz1mdXhgJf1FQAn6Kn7TirsudP0V8DqVV5hyfMNUU/S2cxVyxZ26H1MwJLJIEUqHT9NV
uJAAKpZU6ekVdQNfV7rN3rooszRrNmdnLn8AWIPfHRwlcudn9NtcxzB78QfOWUG+xT5x7JTLF3jv
Mvf5F49Vr5cwgxBZ2fVaYj/vu/t2L2wNWemmwRPI70qeA9bV7nO/7oe6pejkCSk/luhDRAEPsET6
I+tzDTFdvKwMSee8zfIY3uqMRo6ens8l3rmGkxTn2G/r7Qi9bEgB23NpIkOA+hIllXQJBY4hbCN8
5OZ+wWyQdNTA5AiOL30l1bJZsxOGy9szuwrIZqELNQn1KkJ/U6Bynr82Yq7Qtm7XPG4EYMdNj90B
4x+fJX7di8jb/8FxfgYCXa7MwJPEnQKiKkdb1RQ+CcrgAn1gihyEWDtGFirQqkHtNNkfuPFm3j2K
FkjV1FgqiMtkffD36KF6cJ7XJkIjFW3Zyvy+oQL2ap+eC5d/Ef0XOJpI6lrXFZUJM10jfSXwNeQO
DTh5vvFrcqMZ9jgWN0CFzhfrVX5a/yq1KzCTAp7TmD+vxcsyMVekLDQzFO8gDjml6HCWOmP3pLig
ekzYygHh8Fx17vNTlCEnEuDXMonOIcA3FMB3Z1mqlOsM99gGdPfNMP94rQlN7yv+vTskgaXZkZKa
cR9oddrX6CmgKYBq0PuERxntL2wanwzzTFy9WLMFZpwIudt74bRRG1XckA5HqFun0oKJeGsQWFYb
vCM2/PRLeAmhVYLgpkkEEgVAPFKkg9RJ+Sl8KMdE3hJseY5ZRzp374a8d6eyUEK9hYw6kFQFaY/d
Es6EBRLjXF52h+i7u8iak5+adFd4Wpb7xjlfuvszSlwnATsGaqwH/gk3W2TJhp2dg1hAAWBH2HUi
eTbpYCPMBCvgQEf5CVjwxTawpcBLh0bHlw05/J0XvxOW+luaPws2fFZHCpnNpNhEAEjO6EwOuogH
jwG7WxWOSI+03jIfG7gZqk4eOb+QjYau0wDMbQYE0X9kTkSvkgOXGG2cvCyIHSS033frSHmLKf4h
oTGITvFORJasdUID61erPIx80Jerx9mipoO2gWxWs7p1+GHOKYIdJKTy2y53S0uusp88OGPU72Xl
tfAXzK4qnAyUAcznWU5D8XSMQoC3aAgxjlfVN1JZcFiQBTGuyk6v0VbFa8iGv/hOXT+clUx4gf+u
MOD2ijpJa6sxoXiHLqndhHDR0anxfolL0fir4I6THt0lrjSvdY1RfEdbGFZHo5Qfmg/oNMmC3lnR
gkZ5a9G1m07MbHqIFUysRR3g9Ifhi1pWeMvEpNLAvTdciUNw3q08xG0HudRHVigocNv4aOQZ8r5P
3kYudVsLxQ+tEYrBafkOMFIkCaTOZRwiayYr4SoOhZh081pndLxpFzwsUB0GQ4ZiFFuW3Bf+PNC8
6hkqkdc0WnG5YLiqV3dxOZ3H8+Yxi6bLsfdHRqkXH59yD0O0kflxxUgRDXsEKzaxyH+OJizNc4Co
FjPSWzW/ndJlC9MkezH9ezhobcSwJvV4YoBZB0NETg8VRl/+CrOkktHt46YNjkbxk3WB7NgEiUCK
9iRuWTTINotIwqReDoN4UG7gmFEItElAR1dyMW0QXvLgQmVoxY+IGL1w7NrAGjvbR0VIohJMlB5l
aD2GB2EQijg6hjZWQ7EJgdcvu6fX1D8VJh8KoftGAYa9Yb1FoXc+hVk9w6qHx86UkdAjL+LzHwIm
vNYcTDMLg1JNX92AYmFlXjzVw77kUdsy7971Xc+tipsZRBlrGPI7WozKm0Vkz0sTB0kvooZXOtrp
Umx2n5L89d+dT7O0Ngr3Jlrh4xk/v4h6mC+a4RgLVhdQc4RMz0+BYPhWLz5DK1I+J4rY/c77N1Rj
XPPNGHg80T1puQER2386wC8Tpzj10rZ2PsiMZZfAyxU7VfZ2rOAlptX6NGZGyuYA27jmtcOsewEy
IyTjslCvnWO3tVzOpwAbb/yRdqat+KU9jyktf1NYRsAWTAKp+cgjRxUNiUFteaWrvznLvVZK3K5I
UEHGL1kpjgEUs0TxuZ96SAhgk/qJcieYGz6pIfTO3KYg89EUriNAFcIiQC/yLyaPXZtoGdEUAxCk
0zsgzlawon+qEU7Ak9Q6EnJQKuaDeE8nXZRY8lAzID7UDa1FLyo54BA3eNRZ608H+pDfT2xUd86m
42JxCkUCsSgqFlISP6KuPnKLjRvFhmil+XQxTvPBy5CPEVKhVvt0f0Ziqf02g+yXSD017qgpKd0+
0GSzCDOUnGQJq2aIXb2L7oWQbk0s+OO9IsX29eHJimJXp6/btHMJHzgyyYqBrbS8ZUUW/OryrBQe
bkUN746Fx4emN4/5ipikd8qjH7rSqzisndAQaSjfgUph3wqulVPHiAZy96OhRV4AxJm8mitEUsqj
I3qG4sHCh4KJOKRSpZbqeoneEAYYZwEVvUMTceXR9hoj9X9Y3o1bqKrxy9X7MFfHJInSd3PpEQrz
iRKshVA6GzeURUoNGAg332CHEeqFCEyObXSiuSrqb+r59cgzCcWaKhEIE6O3WHwrvxIo6ix/tbdj
L+7afNFSZR42gtkc0/XchjqBBIrPbgJW977iZFmb+BGNxLywXSs2FKET4lok3bDKgwmZjgCcTrUE
hKBk1eTanxNbKQkJyYd+Ou0uKfbXOXLLrmSPlodup6n0YL4J35BxDIZz5KT7aL3RbH5OgHDitMMG
IoLBfw/x0XIvm9BVDQKyWgE6NllscHby3/6l4fKt4lX0U1WzaWR4yiLepL5fh2UR26UFtgtPslaN
8E5PYlY1LSQPZbTr3db8maRdlTkWADL0B+dcLFVCTuOZotlCaXYdPsZL8EyXfihDz1ObF37ramz/
C2KgHR4EQsC1YO8d009dP3zHM7Hf0DPMAsdKlQEUN5vcxSEpX1qvnUVGkjEhTqkZKI3FDwn3XlJt
8s8M42kVJok3y4mYCiXCavDS7NvgBkE9tV08iLRbktH6B88Osri2jEtQpjwbybV0JLWGwFfTpcQr
Gnnd4RcyB9NcW9lkhealIxjGpviq5JVYNkvh/56CqCIfRMEYxgYQoC6rEjxRCQhxI/tCDVP13JWr
GIypUQSXe2h7m6xtRYq/x8p+9GH2Ue+3CWrKd+teUuWMoS/ejN7Ho2Gpd27EXizydnI+HjnakvVx
5wCAL/r/bojHkM2JwG+m4ipZ7tcU6UW9gocIGjvZ4tVjO5I0xnjt+9zzoBaT0DV698jtT9J9MPfk
qFAduZe8GskjgN6hDbZpHjA7JZLOFp2Xn2h/PFQH0w/okt2C3/AVR7savUFpSuXDmULh2Z9WlwtN
sldNiNTUME5Tf2r4HnBh75kNaSNkwwa6MHCJu9wUghl54y6KUpnhhISJYSo+sHMYa8OxVQyu2S9I
vq9Z2ImedBJ8aOVzm62z0Ogj64gCukQ4G5TT1zRbtmY7B/PvHMHbu1hJIsWnLk4kNZIRYCsa4ZOt
bZZ5pQ2dLXKl8WwFeGzYy4nfsPEs0QeehL8W+QZT5Nlt0mQM8kz0spza/qQ6QBdMnB7BwzGjjJpX
gMGApcKt/V2HTIL6Ki5aMxh+SEZNjeU58sH7WuRqlaY2MJgaEVf+7CcW7s5APnpGGwvBmKQHz9Je
5szH2/6HBuf/dS8dJtje6SJ92L6d18+oucii9z+5jmNSUw+p1vMbst7z7RFU+i6Woj+CtvKZLgCD
SHZgyKJGb1ywSKbci13kR88PjVNCt5B0JHE3XpF8LnkcMgulXOmElC18jTwUz4/HbPXR9q/qHnpK
x4jMs6/B25RF4BFuGZsE4oO1dYsPhfhpEYSPaLL0MwyE7MGZ7bgSgQL/hmS9oITyeor0G64SjglW
GrTd9FcWXxQ0ioe2TCAqR7qGHnET3gjI6KCH4pAPyh1j681OC1y+JYoYjoHYA2U1orMPZglIsGVI
+WydtIrJ1V6Qp8KDYLxcvNNKFjwkGzsgJSr82RAsyVlRWkeLsuNpz4L4uinOYZHfdoA31o+zE3UD
J1GnMjjywajA47UqPqxzNHPTLI/OM5HeQcKog+ceGofaNssGzaQh2C+FlJc3fkqpzg6g5F8TtM9F
4qoAtc6+mDEWK2s65vFymAfirHTzn3yKTCv4J4TyBsJMLbwtc27eOu8UtAEx2kRXoIrCcZKR+F+d
jQKd8enj9vKRuB7d3f0ljdqYyXHVDjVPWfbh8wnUEkvtXWsZGNeQ6q7L+AW1AtyfV8FOOcaRWqxA
M4C+geFicmo78AHYATumOPduqr3BfBjz6mnHhqUUqw2DULlJVb3RAWmUrI6vveQ5WGlwbTE7xX6k
tJkizY0WL4+uIcE8uAN4n8xt/021PPz/cuI3GSTbTbHfAmqgUAwdVFKfyygsm1/t65n2FoJli3dV
pjopa6G1AQiPpk168XCilqgUriOv5OwzbB4dg+MzKkayzIGkjh6Fls17gjDcOHp/156vnPZMT5W8
ccSksQSRUuLMrhuy7zhzXSB5GeWe55+XbEeB4CktCL2YePsgsHPJEEMeEKCj1KdQvFNGodp3rIKQ
d3PPgudc03U0sdWBhpXy6vdDBMkyKjsYrufElwYVN9qzd0/zlKh46u/ORo7XOoz+6oZfeXa+IzMu
cH+HV/HOCzwtIBtflQV6FGu+/SUMvOE546B6FtMO/lt3WF+Hc//5LFzbXoYsR4iz8WK9E3pWTTwb
ECeguybR4gsYOkqlrWmV8n6CJN5gMcJkF7qvlWcQuVHogPV0uqJQjj6nLu1gIF8YBpxJ+EL1mdlR
G/RhjUjxYGsD+VSXKta/YYy6FVZaVKz4j2EUoFyZonQOVFy9npQif/pFN6m/dYfyRsK7tSj4nC/F
NCFD1L75vOR82U/GO/mJBZiMGkgcq0coYwS7GRh93tPKdHxnS5aRUEUR2lR39YoryT2uVRpw5ArB
3zMFXDrXjLzwepQWuLhHqewZ10Lq4ZhgJjJ3O6DeWLoYRIHclvS3EYQ0DQmSfuSPcxpHtASGUSQg
KgSszfwQPmpE4WqZ7Q/mGpc+QqZpwm2bp4NvwYGVeeNfB7ZN6IYl0Ioj1H4hIy8DOwd65ez/CIh1
sVCp8IC0iE/nB1uiPU4vZ4SqGO0X6b+kDev1XZBYrziKCU/OaZ1G/cZW0SGxwyUkTj2M6nXlo07T
KXqsjZ3BNwApKqaU/Fb+E6UrrFWAKh5fbh9UEHc+oamOOku9q7bn7otJcYjal5Asac/NsUZNawh+
fjU3nDGCr5BufixJrP8fZtwc9tn/BwVTOoO+mpwPZmzc7pMZrtA0FCTeEKIObUY/dXGy7OwQoJ03
LqbQd9RHyI8BGNQKM1Vqn40IVNcoDEcPVcNrxXtOxgZ8/rMnhoqCAw/+R5JmXkmvMIgLG3cJRINO
ibAjK8p8ArHdMQTgubEio9Ggkhs5eu0x52gpdHBmEDz9HsLm2cHhLGuz3MK3uDeC/eK7zw2q82FX
GwXNEaf/odSpbSRxacDLBz8ioDJqtEFR4ZureDaJE7G2Lw5Lx/DmSKFKu8pJeuXvHa3LdRxgBXMv
m+wdPRqmW0klqLPKvJaEZbPdhLm4dz1RX85tKRbTEGHGwIVY4yb//yjPz/dc/OwHKELXxQ8hAe0+
eMlddjd0nd+gCOrHx8LHTPKqOHcoIcQP6XP7AA3yT73FLomRfnrDLPUOAv8KbGUHZ/MZe+dZeouG
oYc3DBqCzgxvObbIkcm75EU4ZPKgZ/lD1Jrf59uRf1HbOAx9Mip2Mwqijixzd6TtwUQwGTysvwJw
xOoZJk4WZKOTTqH0SsxEbJ9CFWwp1/u+2y1KGyxtB/SDN/vfqwXc95s6VNtP45rWSoKSTQae0BHc
m5nXzQ3x/Z+OqfZPXrmGTaELnARVbNVChDIe9olXJgf/fidQ2PZ3tgiHdlGx+AE3ZE9uLiSLA1HF
SLa+fBKLk+j4RKM02+ffu1zbqDTMoDCjpOrD8ci9NddGea14RKwA0WTeWH7dFinj01NStb1+M8Ah
g2Ho7X16ssRh6cf1ZgXhPg7XSUFONOijn2rTR2sExqZbyGlKmvkX2eNoBW3qbgy5t6rJXMuATbO3
8hEa6n9lOLBrzxwuOxg1SF+TI4Egmfgn34te8jCMjF+qPNYXaZkFPuAcochfaO25OclEaB2fz3bR
r0Rh35PGmAHzEjgojifuvoP3h0X9CHWiNunHzHuAGWU9A+ybhV3//GE3McW6qQmSZq43L8Ac13O3
T7pLJ8jFEGpzMTWcEzM/hhqlYgSeMRmE+/kSucR7vCbeCJS84eLV0aaxw5QLZo20hLYa0c+9VKXT
bOrVHm37aBpEk8CejpN/CNyJW7Ys0yRfqCVZB2DlIH77OoaXl4M949wM1LM6mb1q9v7qf/vYOxHd
wPtxChgLmons+vzKwZF9iUof0UlqxI6MWmmkjMPFN8++cxyAilaTCpbkQ6yDCideNES2602djJLl
hctm9pUDa8tsgKV9WRMjZrWZIhNvKPSTl/iK6JAZ+KkGYsbHeetVvQD8BXaDlt51BOvu7WEUfXpe
NbADtrdAjiPuLBVW/qrBPJbTODWiHGDdU5X/F3A08RH/pFVVz/8hXKfj5lnqvHnMX+yYBzwqhLih
wuNZF0v+wk+8pWyr4c7UKfbJlaMjs05PWBEbQ4zlRIXC4gwWCk12x0GIlbuCd+GWLZvZC1AaG7uh
S2yEBFUlovKnHU9DiaqK+Y612HKW/MxbUBy95/tM1HMcl3O6l1q+5pdJEWceUYUUak4gbgziYata
j5w4Eo5TbF4usNP3+XDP0aRbmWZjndwDYpaloSGEQnFVSMvDnJpUXTwVnwvCAjyC8VrOOo/wj7qD
byb2y2DkdHHojBioCMSRrBXQiycOD3cyh0N2WqKLOVDh0kJUQ7HjdfHBSsjEwf9seTnlXuAJdEIW
++y/4L8qI9EPq0bMNQENJTX8HN6hm92KF2dWpstBDPlPWj+DLAfZKqeiqf3ukM4TWTguGdIpe1hU
MvqYWJSiN4uNNr09FyHCEBIZSh8xqh6fSDZeQuQE3812nUyNPVWdTyOHzm80pEtAesq8f1AG0Udf
CmTtQ5OvlzBCMaGcjLTLAxYnsQ9SPrXrVQFiUaAGgxJwUilE+0SGlt/WayBYe06QdUwf34T2pcMa
zne43viTac+N92niuH8r/spth5nd6HhzKC9O12F5Dju6l1RunBDeO4ngPY6yWXaGhkKQHDu2YiY/
5NJz/QMzs3DKkwrSUjmNroppBK85+LIKCHG8jCwrh8Nz8R4AwS43V8A1/Rt1jJ27QPOxnaG+FTGu
/nob8qa/PITnbMoMCLjxfM8S0+djjBVBsOxZZMxE+FzDbMMpGzNuKM3JkULz+ktBUXjMP4GMyTgB
zFLJJU6mCuQgKdtiNzVsRu4K3rwhs9dms6X1sOXy4PuqcXxwURrPI4iMh95+0Jj6ixykg5vgRpzS
uh1f47UbZLXrNoxAMXkZjba+1Z+U+RjPsPIq/cHxeYzAo4tA/9tUS+n6QHFujXVFCndLi66p3tJs
R/wPPY8EqMBOqKtgTXABelpH8TAZNBDytCJ0b22HsILs0j/usxK0YQZVA2sRvCG5LEvyGVNALZTo
uVaEuADZD4FhvHqfx2Mv2gwN/HnZ16pvLQggAMSq6nTVwr6pgj3/BvdoYHbhynVTwyHubei51iwJ
RjuJUdk9dkTyTF6lsM2z2y5Rtb49YrOi+NsGoMv0JRq4Ql5GsesKuFyc48E+8+AaeepEel/DFX4z
fcEUT8tbYvebnFiCcay+h76P/lcwOdu27kWApRGBJjVBEO6+5VH7MKoKlJQezXD5nqhsv4OLZO9U
5kP9xzdnA9kYN5eFOHdjzDFTyXumxVsfSG2FYPFqIMdjYKHGBBOnUbINDoEz2xyLGTFRNj9AkhT/
bbpWoCgQYvW7gz9ZeBl203IVb21tPWSavXmeSntcxFIHly9fuD3oijRFiP4UR2XBX3Fwjxf6TfVk
UBIKeChOl35Me6uJk7XZhlf0fYRJ4EtKeBrsjNsHV364Jl3FHPlH5aP4uRovR7qoVwz1LUXY661b
HnYh7X0+FoHcnkkLlNRVCKIssuV/AmIuKzHACD49NbpZWklZPQmRs9RDexuuYkeQKz7pAz+ACTu7
XOsnJE3Y3wIs3l2f9xI7ojFROy0eLXnoScE0zp+PA40IQssoLhDO0Zek3avI6ZHHcDFNBzVRQ7hX
Ol7PZA8Qvur70kg9GjA+qxQ7yAWMD4V6EmrzN+l7t9Yqutl4MYQMuruwQh22ekC0uIj3kcerxPam
mfNlMuJmxujpodvdDR1zczx1Vl5uc6tPoMRdod3Gkaq7neWbMaf9jlGCAyM32tDGSldvEXbcs6E9
IC+S3+KYd48k295img71SYYAMPMVnxaqJVdx7mtJdiC3+BW5SkVVGd1VxLLlJNYnhRYqrSBPLKhR
epBp60XrFzC6CTpbOtiHKLfaveDnVwXffhQIPmY2ihgmKAXOHXX9Pffbey6/7op01DiDHCS+Jrsi
HyuJr10Br1VsyvF0xGrYQt1GiKxjEqrAxxkPhKwyuuin/JcI7P6cP/bEavEn5AdERzw0iWEzns0h
HzzCfoN7Y0B6NknOD5SqoqVOk8QKIQY5l55q+PL5BPWvZKpTXi+aNTo7P77SaQfWf/ZQnvUB2b6R
+7l44LF6i1dfJN6rQYADR6h7ibfJpH+JznSEww2fJyLnHpDZAHL+Fg1EyeTxHVJIV/surCIppzI5
Mdv+sOh7+T/foqDrFtrhfEErRpKdsdpoAUkBFk9z6jjkzoVqEZhGWO/AVLOButuVfQnOeA46I90x
kQJcwcaEKHfqTgCSKj3ePOUvtoH72S0Axjf+SQP3jaz6zDDKKGYT3GQSmD8PfHpQokJbRqWwSepq
Dr3URMGXUsoOVKm9tr3BlouEs/rHIkVWq+TK/pCcC+KT9iUk2uABH+9C/vZK3QyVvXYvAhBjK07a
xDqnNKZR9DveDhHaUpOTuG/fvObOD2aMlOT8F71gfk7++LL0gx0xS61n1cj18pBZ/DLNJlqL+fc5
Icg72rwcztXc5LAqIJfCUNAvRELSGuo8NIxZcUO6YuDCF3cj+SV0CeIB0PwLNIaYey2pm+7JYhD7
Y8OGQDVT2wI0K+9vTVaT83AlMprKHGb0tRvtR+YVqTP9tADqQBJ7sdxmg2x7+IM8i3fIxSjE66WP
Pyvi6XTTvdjoygbll2VrIfEfmTwQGNlLE9UXbkJ+s31SPYR7XT3rETLpCP+ajudveqlEyWF1y6oH
lL8qIeDm0A18iwSISJSjBGNJCma3ULRloszDs0Tlj+fX0d55ud7HE6XBtcvl+E8rY8E+n9uIdO4v
BbClCv1d9zQfGbklntK6N2qs+EiQFogx3cHUuLEmcS9y8bygZWWGV5MhBKYIVjL6YZ7MNbH1mL33
QYmV6rLyPHVPOXU3Rqd1XSBT3cBbxKzzRBdio2YSFShyIsYsLCZqqSZxfBgou/65rljOOhm+d81E
f2M1o8FyRrUMyEwK9hQt9ajuegUUC5Z51slfqBDY3ZVeR1GsceKj9hIZrj4nf+UnrmGxps2MhpT5
T1j7NcAI+KMqJk3fbwQjbKezsMFx2Gjx2zIXGsM20ARds5Ubi6YbVL0PsKtRAg/VudZDOuyixIfU
5QTtVQuSjSzVSfVe9Zx5GJMmDbPcB8x1lU2okXC4DEdI8NENLK2r3umOkj39zu0ewB1+SXjVqVan
B7V9aR0bbq8MqSNrghnsPTBM4ocBz6mQY/dV0nb4pTXsZ/iHruKx09H5GLus5N0r4Flz8esFgzLH
JGaKs1zp1OINMZUXCFaYKCuyyG4+yA4/KsUC+cmiqb5AKlUoG+TA7J9oQupEC4J9qpvRByl+aOOP
6sj+6F+HRaGpPjh6DjS2ClZrgqXNMMVVoBGpFql5EN45mS6qPv3gK1IikA6iCDGBinex5dDXx8J2
0C+EbP+tvtha60NaRutlLLd9RKH9AFvmjpTEVjEzGdPeAuULtUiRCiVvTjSRYBTHYOdW3Pfh01bb
EWidCK/4vuuO3DJMRJuqQDrNLugr2AcofZXvC2yzMBuiPPqz/Encm2epXu4ehk+DmNRoNhd5J/a/
YS/ljX36jOUh/gzhMAhPL5kjRCrzDH7XkjVW1qvWnTXp2ke2UCseP+9mPHuIMgeVq77P1kD8/fAZ
bjRYUWXisdNMFenQFGTKgnUV0w86HxOxh3cZy+ava+YyHSuC/lVyqDHb4bhb2RWpJFzABhE/+vJU
ybD5XYVypE5eLk5v90EizTpuqsiA3+hb2+nh0vcG2g626jw9LKhN8VsHVFbODWWEl735UQpAMlxS
5eIqmE8A/PXb5UEyWyaZHugspDUCKTVQCOQtAu9S7cysIfonb1d2vgp8FWO9CkWptdbMzI7BHRbX
6nFyn3HtLdHdpJS9RQMtz7EOzBtCBmUrVq46yoRATKLDcyGeUB2YYCn7UHgXdcGrYJWf7bJgTlbc
qDSpuXc0j8hhnt2Q3gu4PbhHmYM+5zm5agSNeujtJ/RO0WNWwUyGr5/SRwTz0v1vOQinHupQE+0E
1uViyjjISvliBvXINbI8Xk9QTEEhSDI50F7f0r/Sj0tGc8BCZZm8H7q95rPrEnA30RQb3ERO/npY
XzoOG1pppK5DMTXBQRtdyQg9OYgMYh7UdU1WsLfH0n9b0aHDMUCnvHLCRE0oV5U1GxTnY5VkcXPs
aYc1hTtcdWJ+6+HsFxdbyCoQy8eztxdDy6AC1bWw98Rq0JNaHODgRywxufje0ObNUG62kUI83brf
Oyy0ggUF5V8us9eJEHqvFZ0Z5kUbi1HNfk/HGcms930tE2KNoLupnWMkFpd0x9jIa8EUgQjCbcDb
CXdr+OWL5DTgII1nC+NbzvCQ/BsdZroHLIXzuiDJGhtf7nvDJ/SdPG1VdCreC3/XMwVyDm0c9cps
EUoOVhFGUegD/LhVE3scaTsm+JuCd+unZjmf2V/l3j6JMuB6HALQW7nidprYDWtesp+7V3XBeqkp
ZB2xMLZoeqFJp8CpcxeV+JoG9PnZyRtGJSPsL6ym9nWfvCl0V29GOUPxNzHBU2sOi9PDMxcBBmqF
7MzhJwP7MIPTg9RNejDf79pOrks/94dwZGiYS+gkKSDIqr1/6EVLuQtKEBiUbxVFw4ddozd6HXIX
fDA95BMekt6zh4OqEqbCpANRxl9y5kcRq1oVs3E4ntEDKXBsGpczH4gfN0AIQMbmentd8F0XjNLC
6YcD5ig6fZpfnRdPk4m+qtLh2bZWmKwfSMp3Ch/PYVbe+weWBk75ltYjvQAV20izZJr7KUjKdjI1
mw2IYp03/aNnxrSAnSwe2gSg0Ot6vEw5uIKaNFRyRCvjlkZBf/6CozdMyp0mbzrE3O+u2zqT5N+S
d80SV1qDaUA3DxV83Csut/UlnHB3Pp+xvlLHLqpIz9LfUO6dGMPuhcUJSz8muQnzMu/yzjeZwCxp
3vmtAuFgqOMORQTExULDeK6/6mWuRjxWjxXeQsFfsxN1xiQgUt1OXz8okjER1Fw/5MS3ZxbTYt/q
JM+45ouHkBKeLCxSKizXHY0K6NFZispYBJVSORN3y0AAaZhgCTXFUE0q0AisAbIHvphVBgVTUqp6
2mxV54nEzLoXW/VoCk8fiqVMTEfAiDZ1Qw1YAxIG0rJje91rRBPYnf0Dg673QZxs4yhfMhbnQLhU
OxImQdnWizPe3L9rgTlOllQf+RAiRVRvzkW7pftb9cY3WRWfvW03NML3E/f6oEDdnL3K4yTGDTWP
gl5xVfZzs0SNndacoMDEDLcN/EMZGi+Qqmj0CczcOgxPW41fybsiuqCKgVo+i3jpb34wmqi/ioB5
eAgq0CWI4Mo8tURWMiO6Hm9ojXJcH66xgsrJCV1dARc1Q/ijFEkL4XnGczzm2L+HnTJy1w5zkCXR
LrWazc2BZrKwBJsB8ewC3HD+MG2ZL+8ssH+X02tfMru9sBu5UhVGoYPvFzSHZXW23yjudYU7Yubc
SGdvGhy05ogHRcV7DNtBbmw/VXadfxrsVOdoIqIednoFMET64+rddO5Y60oz6COTAHdpNfV11wRX
g3qZghzFxpkCxtKCNpYcQGQ8b0EdBGEE1LqxLOg6dwXpq8OPKmZ6GEDA/kt0FPtq7JPKoVdAeiC1
iwVkFuKSWfCMIxleNR4AqE9U/rDW4MMtoubj6h4A5b1hD5cC9wud9X7ivNvk1j+pA1r7Tpj7Qri5
HqJK1gfMokoeZV4Wl+4PvLF9bRD0Mg3be2u8AQdWUVLPRtzlKdM7W+jzOzZkzIjADzxjTnB5Pk5H
4IY6EfzVC/FBL4c854HH4JEKgGt76ZHxJb+K5RSiXDAnnGf1nlNMWEfiYvv9iOM5Rso294AXq+Sr
bRPd5y5ULaAQDEinWcZ8/EWSThZIzMhQ3lNiaBm0nTy3V6Ci4YLUT/Vu4QkK065BY+HSy1RHfUPE
oNfcOI5L1eXS70jj/wyRen9SVwpusXy4ZpAXJvCf8kslqLcTbKFwTSWm1s831XZetIPCreTJc8wD
eQAeQ7hCWrZDMZ39oxQy5hnVlb5MIfzhochQ2bTGXcnRSNYkF6va5eOgmrejA/eqZP+ICw1fYvt+
14z5rRx7p6/FE0Qa+87lqRPUd7P5c2R3Tk9YqSmlGZzbtxx3EBdx2a0t5Td0l8HEKb2M8AyMaXqj
D5fBsJwkbvun+K6512v1nFSXYfg2zaNBOwBfOhqz3y/4uBYgWWOzr/vDo7imCzwFcUe6Xm2N8cAB
wF0vaJB9QGcUtxObYNYG+jNOcHJM8wCh0S8n3ZqT9MwpyQKCNMfvbMa1eCa8astdqRiRZlioymbL
B5lwvd5IA/YFN+b0IZYTPUxxOUdkSol8MYrlRTLgN+Lxradse6FEO/GK/WW51+zMS8uvpVtQuMaR
zO+CgyfUccbMiK58YD0LKEAUcIUq/LZ3wTbLcwHwVG7pktrJAS0fNzYpljPIfK+dle/l8iqZpDIq
g+b42IJIret54JkU57+hWMbFFgYg67Ucuth0hHIvvwIHEcw2aoSpmtmY+xtGBwwQGB/ZBgJfVuhx
r2cQfp3AxWt0273xhldoBkcC+sE1UdLA7HlmU2s9jMkPFnKXtRjo3RCySPlWEhPTjrEraovKkYLc
SSMuaZ4m4zBdHZRUcgYNArpeK/wqMsvemTEKpzgMYJGfXVnHiSTEfmCb6ShqNuP/zOLwROsBekGL
uhLOPZNLROrZ8a0eDSjygJcyCpTiE8Y8ZxWKxMXCuXeqV2++D9ooRYLcI9zOtRbnf2/waAbEa/8e
uLmg873Sw8p7d20bEwunVPNn9rJwsi5Yi4sUMB5UdP1W2bFqhgErYjrgPdckk22JQQ5zaY9SJ1HB
0AbjrWhTUqyjMNzq+a9VLx5Vm4qaihuhSW11DGnnkIQbekFLA34SpUUXRtR90N9HFfUlC87V+A+V
s7e8WYWyRYDawFReJARjQ1SsMc6wZrlj3Jp9/AtLLoWtbtV/lquuo5Kg+PZiidbjj8/iBrj/meLZ
M+1hmaX0cC3AeN/Jiy6zNwVV3ZuWfepKb5Zy/CC3ii4RIb31X1cfSvo+8HHHjG67qJO3t6VCuawu
z/dsiu+OeQbpUy+YlY8gVH6UtbvgPloojnNBcJjSd2UWGShL47RDlnzbnb66jeeZXmoW4Wrqe2R+
SEKleOnFm0Dm7P7HOUW7WthWGrPHni+/2sVIGjeQsGPPrB6UnXhHapb6l/cVrGRXBQYIl4Q8NhP/
fttZohlTahilZZB5KkdefT8u/5Q5ADyV8PAaDe3JiLKDvi9mzWmM2Y947QHha1UPcl9U2S8UCsXm
tDaYdvRZ1jmdLs4Z2OIAU1BLgW1pW04ERkoEqkTvnTcdSWhzy2sEn1/M87vo2u/kX+2+1j/4YS/q
bn89UopjXebUP2H14QLm5PJADo1ljqGKV8/RjqffyXVGXhrPMTywc3Ws2zlkjUXtEmMorox7pVcU
uN1Fk8LCoE0ioGUy80EG8fVQi7GnY02jw12izODQB+bqXCuncVNU8CvzG+iQTVhtdzxvS6zRWFx5
Fkv2cu8Md6rfdbWH9EXyIxFeD3Ku+p/H1MrZCl/Xkz3RCIr1DbmS56nj7vbj4A2iw/O09LoHR04M
xwhB7IbFOylTYaMhmH8EP7XjNUtsPixpDNOyZo+8tq0JG1Z9UXgvCG2FZ8alIYfvAsC4tudkE/hM
8j6OZ18dk0gQHstz5PRdM+BrID1foC9Kn737imU9h/Ot1SGXKWc3msrUcz4/rRrFTmSJn9XvzeQV
9Tawy/RyCnNt8Vb2Bk5qMon1gAhHUlGluanYmdRX17TB13vevv74/q/jbfSoNVz7RLI1jyVlQqd3
oNX/0e61Fl5ZVO1a4HR/eXUPwvBI9LaOaR+DI1novbzNIAKpDC/XuTGtJSPmjf/pNAZrEoggy8Jy
QtocZEdufBjdqwNjZZQloX49VljGMU3Don5Iv8m4YvG83FckDZtHpQtwocvTDe/Kc095NypZTgUI
g/p9+34E2TebZzUbfUL2aOHmP5x1yMpPxopC1KvgzVhDU3pj7WRRgrl1Ghp/xLoQj3CMfOPU7oGp
59qql5BzbRdNFaPpu33dNktXW7pK4nWGGh+gpAa1cryDkLJrQ40VdVCVw+p3QtNMwmmoz8XyWcHJ
doCUxle0DgNHCabOCyILvulm8qDDCtWsML+sqrkFCk3fLynPndaryaXT3gPm7Te1eRoe9IPcWFUg
q3p029onhTQJ/ju1aH0KfKbag1OHWWRJOPP+dMiqf/iKrqsar+AmDxBEZshN/+RO/pHIKj9pDRtR
/oQLtv89Bpd44iTrMuk2yy5ZseWl1v5/ABO1/zJLOw2Y9iDDawwb752mQMFXbwl2x56TqnLO+Wf9
EdJz8jY1s6K6MILySzd9cFXa+ipgZVxdd+5t+C71maJ3IbZoiBMml4ZYdGl7Oaq2OUNDmPIQONGe
5zjgH9m6lT+n3MKg3/Zj+XMrhiMvcoYMDwT01CHS+MgqXiL7+VIueNtYl/smJzvnNlTnNf+Yz1lr
Yy6fpBegaKHHfrRnlGPAVigGOZn06JU+ZIDAC35jYUed/v8h9DGl0l7URvQnntOCRGmND3IuYQvQ
HWcC9XWrxFvT3K4zFG3jowp0X1fFZ9KCc2yF8s6qDVjCUmDoYaIFzga7ZR+/35TO246FVMBqL/Hb
/RBETwiVtQ4/CCeFB4cOfmPMbF4orhlHUs1nwHCBzuBWxpTeebsxCD/tzHfaPrisGUJAGUVL7hsY
9hEQQcd/yhgQUoFbZvkAzr+xrVlflva9LArubn8cSA3RSEIAZyWWfNUzuwICk4APMqnk9woFQnVW
5kNmXNNwy8dE7/ad+iu+5U0lTwMCQtO76cLpvOB3R1VB9qLIV0/0jGUTHKuXZ/y5JVeufdHC6FqG
dSBiScVp7+VI2Vbh72ms0qi/VK4VKVROVVKL+ZDF6by2ni3hnCNnisC+NkjpeHsovUlQp7RJ5cYJ
upTI9Dhpag6m1SR/7ovpZJ9h0CSiaCQEuhfBtefCa7e7yYuRBcIcCOnRbLm1swbD5H3bht2hEwEq
MJG9qY3xZflvBpH5pIv8HMaoXQ/F1A21kOux47eptokvqHmxo8YbIrsbZZ1ymlThBT0qyvM8qmVA
UHuwuBr2q1BcJqAK7OtmvfUOlA9ZNl+pvtbEqIgQNQZdv0tp5bgYsQe2KsdDc8gg71i5FzWflii3
iW6yCjbLlJVXdcL2scHNn5+AuKc/mK5HwHrsuy27pm4OMwkzcDd4/JvP8cK1g3fg7BjxV2zC2b4F
vA8j1HqhqYpNsoKTtA+SgGC6o6vlVEIHKRVeP0AZFJrCkGQpimKjCgI5xF6Vy6g9pavyGC+wVK3T
A40jsl50CVYPhIuW/4b2a+rz8m8CxsO+0nHwy8PHgISPTHxbFY4OivmHj72rIEyInHqZzft2ZPZO
GGfNU0irrOvEWUyH4QlQBTNJr3FrH1HkTmZyF+HyLia7dtBYNbytC8mspu26nYkt6Qkr/y5ej/0Q
Qj8KtS1kGmQU4bpsii0864KBW7k22p5Huk59s/+fmQqJpZjE+tG40QjcqhFhBvAqxWyTNQr6Mdda
X/WotRe5bKN+Q7d6Lfv/7dPFweE1/ZZ8k6SuQUagU38i+dIHdS+mniR118kUT0DhUo+CJZKTOOTT
FiqQMMDUn909331eHLO+cw4NwzCLWEs/f7RL2gsqh1+z4Lmqn7oPuD0yCiXS14ZscB2k/Qbw8dGL
qArFMI2d+ENmGdOdwwdjY8uAeH9yB6GgSdYY3ZWLAt8v8hACei4Mqc1uJT26VRubc0ZCUITclOyx
P7DA2aNwyzuAF5iAOak5OAA9i0nqc1gWPl2jFs0eGUr6lv61byM2Riauct5aATezcljhmg9cYuvg
DG1bSB+SBXH6yE+ssUv0PUdCTAnxxrAGpjR44bYjzQYhi4zhF27y8gzSM0+q3x0AKbNEaGZmT6lS
jXrreNj7hTrzWDG+Ln6ytWs63K2friepnKMe9eo3lAxMLSO0zNYb3AK6kSf+SimtckzO5WBOWs5w
IyG/aJVQ0GINI9Li/TvbyVXnqFQYqeJnuEYRvoT5XgR8e7bGgIJYsCVmOJZ1a4xvUPZSxdiGkfNQ
88AntttiXQt1RKxf7Gm7+detXlOp4gnkVpchFQhMkttkGpfP4YgvKWS5tJqWI1luzqNdhDMvYPec
OLqgOuxdFmV/ARtQPg2+iFmlwmRgyxiM6TRB13InTwJNVOIX2g4Lrj/eu8uQmsNbKS2wDUPbPlTa
+eErNavlqmbCQ3g8UXA0Pvx6z7SDazrgJSDGruZV+haa927FUo9Jk5pm6/HOekfZI1cOAVtdd63F
+LQod9V+AIR4Cc2eiYeoD5w2miGDH6Mdt1DIx3VhHl2+JabroTg/9Zz3N0GXbknZbvGhpxStfLMJ
zV0VDX4Rzonc3kRR8SjuI/X0lqJWaK5dkp7mMr6WNKz4Epp4QZP53bru45X6Yx5hV3YmS6zyRLq6
VoSfdLzZDbFXuzTLWu4jPbB94i1Kmf4A3ifHIYJ73gGzE5A5haX8+6FBNpn19ZcjxTH9I+C9kd9h
hKwoprbgiUjsxmgeTqavbSj/53qyEIg3iuLjXSKXZHQgX2Cc7zRvyncl9ELqKz3+qvRy845i2262
w9Rvq0gpK36sgyI96oh0Urh6t+37ciSDVBbDPiDpNKlgHc1eB0lOovB6IBWJUsry4o9AknL2AuOy
AdyzopzACfA+BWyGsx5DT2o6bkog8UmEhnTpaBaqwp0grig0gRSh2lyFVoFVhngrMvCcvlDNgzc9
aM91NGXY22uvzdmrRWwBUG89A0u7LecZDOjaFNF53XuurNTMMuT4We2hADCWkrT2jwNDicr8xWgh
2jSUf3a2szrhdil0HRX64FY4yyi/lPFvW1KxN1WYFQSHOWrunWyDiXKS26ixzuMvxDBiu+NRjDSa
xECD2cSPM6IJebiXKdekC7fuZGX+XmYyoLSuixvJqL1dwEGaDdW1PQHTr/Zkn4prxSh2BEuRAXKG
SVM2wbHzRY77+KdksY5EYcYxa71hEdSTt0uoGch0DLCRyagG3cPPHXjE7lVNHLOgzD08fL95ELJ4
Ymnyikvj4UosX00gWH5UfK6PuafypxeeIAixTfybiIdcSs1n11nqB7QV8fXnHaahpZex3/8xZlbf
oqFOUeYSxVX3xyo0E0OpqjuRtkb81Gxs4W4AqFcNu41Lokxm1yI57Qabt1xP/tqrZP1KWfPsAnvd
i/tzWCy4OoYKhsr8UDosfjyKAhwsO2IA+zOC0ZeE8a3x3CjATYtR8QTTavCfdxAlknYS472rdzeY
R5xszQhpSs2NSDUo1c/oHjLfZHQL6TiVZx5I8Sf+bKT/3Iob1F2wzlz2qpIsIAfDiZ2EaUgjPBAO
XnE/yH3ZfJmKjUHwR8g33/0Aihf3SyylIbJA2gLxh9DeFiTjrGg3VBao0jKhlKAxcqy/hX8Olvss
pELWl9GfiPnobd8341624wp072FPSupj5M2HBiQLULxt7WXmXCVQVt58BvFfCC5dyzdMmBdYVzvm
5gldbr01Fm67HvmvF1BiXyuI1VJEFapFDyLJmHLAIwR/xDd/vMSLuvv8i93qRck1/xm3g1V0f5FJ
z1rNUdJKDGQLzbCFIbr2PjINhhdlZOqaMhLGXDAgE0OhEMrJv/rRQHPWN+oR7HwjY4NMtnR8MGXZ
1q0LlwAgYJBOz883+veEU+v71FjymvTQFAUR4nb6U8RGruvvs0/WlOlzJtTFBfjDeXLt98vGcuzs
4BEFJ4IgkpAMeDnQhPoHOefk8VcYBfukoLpiysmeXID6rz98vaBLvP02lgkHKU9H8O5KXVDBI99t
T9OwrTtwyWaZVYJpxqJHpniseBVNqMHoQO9W79CEcjPHBzmBK6OKJPJ72fjaB6eFwBPPqCnNY2gH
lDzU3yf80OiPFTm3rL4TVZi/XP6lPMvDJuDTGUOfPzxMaFlQ1z3nQVUkEPILauKw2Z5vL60mbiFK
XrAYc3Ci1W1cI9lzQxE/LVSIKYXAAVt9TG7eIex/iaSiFKvt+ESbG2Ht3mvBpq83YnXpAYfoJa3w
HISmL/2/xq8habaRYkiXJMCIu4KEsIN8EvKvY34zJ+7Asnn/BEbA8tRYzBESGZuPLbDHIhd6oQEQ
YFNd3ljCuBveszQEnFOBeFgMbic+WCJbNPD6XfO5CTLMg2+KNM4+PSk0fZEL6Gn9dMTqOTDd0aB4
VTgiraBhUw6nKzF8bUYtpz6owxLh806yvTp7wjGA66cc99+/yVNWjnXWqcz1cxAZR+fJW76gxzOY
UmaiBpVG65CyU+nYW7KmfBnlGCGzAC1F5L6oKvQtN3MNlcluO8M+Y/gRwp1h1a1B3R2GOA0Cm39t
xTSXWkSLKvj4UliMxOwLq0Yey8MR8QiIx1Kt+cpwNfr86HAQWyPZj73Y8BH9gD5/7rqg/S65MlJw
0pak9PvwvBPFsncBVBL1WPdD7LqrBAPQRSalFffsdJRZb97VaQXvU74II8MrZmUm69dX1yljTcfN
rGGKNs8/ZHGZya6uDVZTxGQeogrXWWk51pfFHBNULwPaTE/i1PjqQS8SpPvekLLg6lrorXJH2Ea+
vHR/2FXUIYZJgsqkiq5CQYBOzNmVrZTIRMGYgwCCVElHGmLhVSDVJApAMmX1cOSIBFa0kf4G7UPU
SV8o7qXwUVch1hLWax68Yro1QnjnfXhiYbGxCNV0N7N42wJu9TJEHnmimdyl15Cykfo40arQihub
thRWP0wALtrjUv1xMy0ucaqmPh3ACOl2OYsgctFbknCH+qRWczD/iBY/fk6MymSZVEaM8OK91d0O
uadnqNjq2fhel5ljqaOrRd72qiKMnOlIAQbIVB1kHyQ3UOhnzlLuYxdeTazsWluVZ1UMeAhL/yys
ztYwBHEESHhcNVwr2Vs7tyAUnDf9aYVFcfMbAkD/PA/m09GoIFrMy/XWSVJVfK+2by5rMBaBSA0W
H1na8jBJ5qGfKr7ETrWqCIyirK6qYFjQBPIBTX8K+8vKvTt7fITA2pBWPAmCs5gtjUXI8Mnzjuqr
oorraBeJ+rBfyetyikCV4NyOZcaF3R7hZ8E6Mo3t2v7KJWQQurirKTtu0zDWTv3wb+ucQ4TqRrHU
nB26j4h1UYHEzIf2lEzoVQrWxNFLYAx6mFIxTOYku9BlcFsdprhBTEjpLpTbZTseptgV8VP6311f
4kwaH4qhyauXFkUaFk2W5ctP17UI4cpKBYfP3aVs+arCyYDDX6dALmVpYUL3niiG7YmcNj0jEw2f
8zxOR0hs0gyAY9FYknJg7WPj1jvH3XsgYYCGnYWIxCwg3Gaqiotq2W+k11SjLy4doBLLpQ/2Uvx6
nKUg/lUF9MZ4wKGq5aQL26HVragiJe2q8ZX7ktyiHoTA/eDd5Y+YbVCW3sw8ueI7uvq/T0Se4r1P
8uhuFlBEznwQ3iwY8ICKvsm0klz3akbnehrRPWgt2zStAfxxLLv1pKxyzpbJ5c7mPdkTCBpKWa9H
gKWin8pHXZcMPegN/A+/HrFtdPjFDCf302qB93h7Lmyh7mHbbZA5Jz/qkUIzN1Av4kznFwrLCVb5
kK8CfT2wYAwCVTkFKfMS5TfBLgnJbi5NLuu9cNpvnTSQqNRs9nYlioROCDk3m9UwveH67pxMq8aC
/LvqEzwR8tFG/N12FALdsTGNCbekvvgQTvYD/J3gNij/YYNQ5jUN8uYzXwROaN008WR5eNfb4e3y
Pt7cbv41PCeP0ngcNLF3Bo8j0FiTODu5EKVltTaF7C7vKIkWKhYEOSjhhOPWQNYmC1LRuSkPeD1D
VMlTtCvGmZHQtRbQ3UeOI4ZprAJ99laPrdx9Z6TiUkc4xPnpC/Ufbr636P+Mvae4PPCcHiDdmPmX
P3Q/OKnjWSneX78e71CLnRouAs1w63lu5mR9yq2QWSg1pd/7Jc6W2K6b6ajQ6SNq4ASiAIkW1QYI
x7mKX7CjXCMbmPEaLasTokSuT68Z8xzFsMtvVztD1qw5CxDmwkvhkCtub2pTm0+qzRtUcqzft/Ib
mp+4me36vwjhTHkfYF8Kw3GgeKpWNculBMT1jbpsyVi+afQ0JhiW0s6y+tJJXmTP4sgprQ6/C3r7
BPJun/5+xnUDO8J5180006HqN0bTP+ruFxD05NnuGLmetze/l97Kz8Pj1vsXFBH9HqdjVo1puO6N
L0p6mZfD4BAfuy48nVCIDm99JiNmTCc7ChYI/6ccFkpim3zasZ5fTTI2VMoTCGQtDyYrCWSLiOqZ
k7cQYYd0Szm20Qwu5GXcEnPTLw07ja/TnvKqxXCTxPR00N2YQ3eQbaU9KC2QxkOnOPedIwwTweZe
u2x/FoKqGjI4weydEtfljVxfq9fcwBoj1z7djCZJXv5r0mLcKxlesLbkBsyFL/8Pf6a9o3zgPy1R
HQD49b21usGQlCspmFayl8BptTWVc6nbRUVJz2ZK/R3ldwW7RjpLDxI3ISo7zO5AohwsL+2MqX8e
nOZavwCTEwzLyMEsiayjPqIRYOxQ3YPrSfcu2abMXOR+5CAfqJr/m4vhiPk/o+EoaQ6SmSWWPX1D
KRnLDLp5YtP0JjKpMPY1Xd6TmV8PfOyC5HlJMBUkYJTH6MXKj0pO1PTL2OyIBydEJUkV/SQZz1ci
0zoJknPEnBHSZ1YWa59kWcGGwBRUdjtEXCw+ztJDhHA7e8Yg5BHT5mB/Fdx2Ph31Y0ZrlmuRTI7O
noHj3RfL/UliEPE/ZC2MBhOumfRTPpyj/Y6jz7iW9vVcjCwoSt/Uec011qJRkg8DEKDrO98kfJWj
fCR3xk/dJIfEuXUhLzLFFucYn8T79e5mCJ+Jdkh3dB35+57vU+m/xT52cFAiEt9Yx2XfxioKfmGo
mtrMqDCI6/+zwGPDEWgxq0FG4gyt/MxG8nc46N9+J/vehqfeG/dddTFEWQDLClu99vaewV9eKMmr
0FmDzq6iN/JenhLB79+tCZuwt70Czeb/IC+00/56aTI7NFognIfWbGuePwVcTPTCaYxTU+E9YZGU
olGmZ+8y7xMY1O2PKd+dnNfh/csbf0EaFFdQ1+mGuxlzx3+m77tffrs9XDl9Jp63euoHCjyL99eA
giRF8temx3opsqfp840YyCu2FCTpgCvU0+9CEMq1NlslMs555prEhMPRVZUDOKW2f6KruI0aO7rn
Wp1GCYpLkqhMC+3HOEg5x+u14v8E17qifA+C4X9IiQRF1a7pLav0rQvpd+fdn1YrhPhcHENs7rVC
CHL2GluCsU3krtXrN0CFmIgwcwe2C7keJkCnc0TKZoKz7rclqc8R0KM200SIqfvpXpTJkkn9enEi
p3YfcqNmt1B+0FYF9FE3c7NNiTq17wvXTu4quFc+7Wru/ypCX28kkn/NN5ntC6YuijoJgjLQdQTh
ptrfgXH1Hc5Eq5xcjCKc1hHc0vqzUzJGwSIH3l+gok2GAOzjdRWBkRkggvOcgg3zSm/zn8/UhSTC
bLHOvUHBYkJ9kwjJfragv88WUrf6a9UA9Jvj0oWGibOBJtlxqJ6DMzJUTGBxEhh7+tI+ueyLZPxL
KP5FtlTdp8RvjM3mTGgSwMt4+dXmgRxe9f2kEu28XYT6xPcWxiUdH1oMVSR/0HgI4CFkTxrvSEEc
Mj2JCa8jVfwfktnxIU73v/MFACNeE69Tp3dHvMxprkHMFCF2j71k0k/NxxrcSviasaFvV8ZGA1YT
mpj3KZi92K5MFjf/AwjgR46423H3iZF1vM8og+kZFVYossrfvgcAwy8DyHcD3M6PHC83blcintlx
yyYWX5IX++Nu+qgHi0PM1tr9NB08FoH4DShUIaD/xl7FiyH7UVpqGyybp047pHc8KyUe7LOvirGZ
S6U1zbTWLxI6Ae8ISr0F+ciNVtXS8A9OwUeqHCsI+deu2M1AflCQU3pCO3nZol7phquIzlVFgRoN
1yfBm30Rjfyt1o8h4xv9o1SJH80aBEOhbNi9tnw5r4yh3Y2PIsD7xUfROTBpNH3Q4EgFyvWu6Pu3
wpOrYlZo0JzQKJIUwTiAKreNxI3J7g2153atsF08Acm/L35NlP83QmblvuUGBvp5rxX1cLl+xxe4
YxbLrp/NFTYv79ibZHstwuTClHyGzLg7rYGmSKDQ12mU2WAsbhALoFKsjwrVCnZqSQMjuV5WNBk4
erNN0pko2EvGTl/mf2hJtgoDKx6vk3enbXTWryXVoq5CPfDNB7W0N0Z0QgIS1PryAI7cBdgizKcg
kWZ2aUNT53sl6CdxqO3vIDYp+uwk2/nLfp3ayRIWRSpmwCzb7+70i0IObZBPB8Q83gNRJ5dgnChV
m756mHeYgx2Y7OzhIl97lr6pX1DJfp0fTtbikZZm62sUyk7f7KCF4g438gGqozv5Y3okO7FNeyUw
aFehKtjw9nImSF1wZTgQ9UocC7GvgdLkwdfLHZzBxnUUEHeMcnYuA8Gb3YzQN5G/kmHMdpGTrJwR
nfYHDSkACITOO6rYNfwRYi2rNRmX0UA0u1zTwy6IRaAUA77QtUgWG58kBWl+toVgl103Iq12H+4K
uWWqrwbUrFgHIW7Hy6++pFS9Y2WshRq9p1xf9Fl9D3vJ4yR9il6Zw9uRwwfvzUgHJ6qsUmdpoyQu
Z5D+yodhJoceH0/TlFPLHaRRf9Y521YXBUS2SlJz2jTgOwBX7eQfzdLg6hhUowFbqhR1LYH2Qeng
Q3lZdjka8DJBeUErN9k5osNg3IGXgLhtKNYgHVJvmxtGz4aGj2dTz2xV7fFyfrIizRb8ioLScc3o
MBLDZdN1oMN2Jp252lDMdRZ3k3W6sCPEatlu2Mkc/PDzuFrqKy24U1836OXophOxHa3kqmD9JhiC
GDfxr0vxXFb0UuubYhREUb1BZRhzze8XyLnQO9m3UCqJln55nJE0uLsj7SPho/CEfkN5wbB5znxU
r727ytlxsVSt870LAD11OKs4UELQPiauC8Myk/96H5LlMi6ASqtFxluWYXyZYkdrLsQC4r6iBWio
9XvHFeAjx0bEK21sPj9L7bwy1iXHRGRTWuCSbE7sHpG+N1zkiyZnJ1qFNMVoJxGKbbWFEqB7GyUX
g1rck8FoQ98sq9bT/ZnJZZTjcRoxIeblAGfCvamkvMVVLCCNCnuKWIgsNMwB/3Oz248cQU0KoQeE
lg6sWVCL7o+JwH0ePyz94VI1u4ZYj4Q0IoPXUrjFRit16o6fLdWMjwaUg7Rbj/9hl33tTQXXynnF
51eWqEpOOK8VvloOJsvrBUo8RpEwDkjw9lyzeL/+9X0Km3RekC41wiEcwByzfpIrlkqpwArgssM1
9MK1oWWM4fdGa7C7JM2p1qAb/1v7Nrna/JCPXA2eGbkN/1/cW5rlxTqJ1ocqI+y0OtKh1d+c4S1u
NVrEPJ5Vcg46ZZC/w/S5Ng7nX1E2yjWcYH6E/gg0nCM6GN1UJUzHZZtmysyJ+Zzf2P1kZA3csuYw
KTRU5npZ4rOeKXI53on620FRtVCnZFNDUIrnt/Ce5BdYovFSoG2FjH6uOMYadaESSWKk9hAemFLe
l6fjroi6lwO+VIJQM1PES1Ct+wL8J1VMLhYKncD8I88PEhI4/OTQ0xesP0Bz2/5c+eWMNoRLA7Hv
LE/j0oiMhCXtEKoeOsZNl0dbVj6R77DjkzW6w88dUyM5zfU+aqvo90htM8e+VJ9LfEyoLM9WtdtD
x4TLmtjryzqeXyj5RR4ixCbeVuUnoyp3+xWzJs2R0lyXwp7AAmduXqdNIfxKHrj6wFgWe9jQVu50
u1RvuhNvtZuBIJM6htrMVz5YLf3hwMGb+DMdrJnURSctY3jHJYaZVXcWwqXzZIQH8bdR94ozO4FL
o+ctdAavqKo88VoAPH9yAijyA8ISG9cl28j3iOoJLW68X65XPoNcVepzy0yBKNsapYSVj/HPz8qF
+Bye/wVYL0IiWFCliEQRMqb4R5xlNXw6IQ5oLLZ16sPyvhFSb14a/vNmg8B1OdAozSTWHl+kJPpF
Q+zkpsi4xr7QqzMta0k7jLQUTlEAcytdxN4dF6lq9Sgn4lVODGDQUM4B3kmwFmk+Yw9qtV5fo7ff
13WI2Cd9sucs/CpXmhnM07yYowH6X4kQWRA3V97K4MLDnxipQdXypjDVUwhv6PWT2yhFeXqtCkpI
X4NfnTd+8ttK+632TZU3c0gwgg4j9iQvAZG4Bsi19najldQVvDe2Q788rgzEXRK6AcMqtMHsYldU
0m5K8j+DFbeFy5iKk5MJrQy3lQmmilfAy0XdZcL7fYv+SK2lFTKvJT3alWs9hel3XZoWPdxPnEsF
swwiTwOu7rPDurHURIs5hO5QZcLtz9wPJod96C3Btv9y1R+Y6e+QdKw2KkzR0dLSkHykydBmWaA5
vFlXaWbXqT/CaeDaccEHOJw1yuiBT6fM6LmCU2m362+6StkzSBEW1ZPH9QHV3dEmXf/5bS/7gX2I
nYpAmXjHfxhMMIbMUYMwpEJZRZc86jI9VRShTW3w/P4uZuECAR/SO+M/ygQZ6/HSyGy3NFohWyff
BVjCIAVPZNi0VXVluolhdKL1+ovITtdnV2VDeTM2XjWlQDCTfX/0P3N8ULc3QUPS2e5g3z3YawJE
Q5366fdvPYeWOO4Ow5guDUl1+O9fdJNZ4s/qrWX69zeeRB2jV96JJQG+ik/QM/SA3AcLVF2lQU54
Xn96WtqXhA5yY17HK6p3fXHV8utdi/ncQQr0vSi00m2jdebx+zVXWfqKCDcwlA7k25w7SCwyRJwP
QcPwYybM3uHuwAy7Cte047s+J8CQc15ugMrigBUkGyS1HUmmQiUfGwh6+uKxAJpuzu0GYreZwiQA
kHR/xO+dateUKhaHZ56L8FtsTQV80y6BiuXowsQL5P+3SNi1jd57GAdetc4RECXloXkl4exZ/Gjk
XvCkPafQq88zVn6ZaGbZyv3oeb3PEvfer/tQAVWvXsJ36ufkKN9dgg81I1oXFTcgrM2lBmpiK6Cy
2BtkXXr1qCeirSBIWp4HZnCscMmkZ2cL/T9Y8NoXl3U4jJupDO2HaDZ9XBslspyTHyncHdMFDSBz
v0k1aQnVz84dqs0896XDJ/bgEMIKZ9rR6SmtKqmZwJrJee6bxDNnpmQmSifdi4X6DyGDY7Iujlfc
aJR1owO7XnH13FRYeMyKu0ZcaMjxxgTLxMbO5YuJsqERcqEHoMGJnne7jPqHUDizC5ByIZ11rxmc
53k3mjeQ5qi7av+KjJVq4YigLBgnDsp+wlhTD2/mOZ/5c/bvrFIqK7iJfaW6c58HdI3Zaur0exG+
aIS2F5ettJA4ckE/wa2+/57PuMpHo7S/RToTGaj5QG4peDiIhnXh4XYZ9QWpG6oc1vhpVdpiGn18
59/jGGHS5HrqFog9qfh3Y4b2R4DZLu7FVvCU3VJ1ehzmbZGG2BUpzmwRUgbhZ4pMKebvmuLX5HDn
L3s8g4Nc/SM4RPKIV2CZZ1q4Ey+QaVyD1C1SR0+5xkUExFHcwKf9/xe0ZDKcfI7h0Knc8rpl8xz1
WsqVLkwCI0Xq3lVjLiGCFnDEbb2TZoj5aZm1MlYOjX6Hc0XKsMZp5YfruVh50QPZXYqvtzz7a927
fe1UwMr4M5QJ5D9uvxJPzBFZP1Tjosge6XJpA2GWklGr8evA5UuxS3U/pEKyS91Fsy2yTca+X9Su
YqXPWz/XvW4NHPlaBXJ7J++4wVeoVXsjdrxwlFfkvzmnicPyV9Pwmyt7cIh8s7ixs46IbF+bBO6L
4MENnAYJkU+yXonZbVmycV8OUjW7/w2kI07DjYTvel3KSh11fy26TCo60DTQbpEYQO7StNpB7RsP
LqKdt7ecs1Ty315qls3yJc/Zfl6wlhcvIZuB6fzDFwfFDju0NuHyYnQY2rGtxU0g0dbOfmnOtDzR
VnfiwXfUMwwv/kKENNpSBhFWfyWy9oKAo2TXwXKgkKVOBFPZaw5FMMdlhcWhuQh+ym7ICFsBwPNv
knn0E3xdppQEdg11Z6Ttm+AoPy4zrtWzcBThAQ1n5+zUewMvmqwBr/RoPFVhyvwty5g4/gJS3WND
ot7anZWHKNBtKB0FhnynolwRGsynlV52o/zT+eRYxYZ7JN9ihMToglv/4nVGwiAiLU6Vp5vd3IzB
FQgNFHvb6BACm3P8fK8Iw++00kUdzcZkLfIJkO3W2fqQs9mgX+9Cuw1U4MT+7ZCIDiyoigGqnYj5
LIdcArk+rgmnguR+NjxBsNtWvp0S+trkiId/kLA9CJvYQP7RW+s5up3OtxgCqsPl9yeuiDBCVVcH
oSYhsZX9YWU/Sq6H53wEx4XexZ3Pf3YHNDTpi21oM7nNcgtLZ0A21ykyBv/angwSMdPjH6xlV0TH
5wqUyikkB5S8jxsZ1uS63qPlzQet0hp39qRJjI9E36GhmwlsXUterRBsHFI5szqT9KjISEZP5nCe
UkXNLcL9OS0znXmykDJJWWOXlRRXMvc9Q7nznerEJLgpaF6SyKaFGgGIfTumZLYwRaMZLcoq9sVC
jIzk113XAcOiZX3cED3djsfmpRPzzIMWUGf99gZy2ABcF7rp9Gk/2g/LlmDaX/LOpGO77hnHDmQg
8hpXT45c6/KeznhS4AV922VFUHXhu51WAARmiqGKIqrCyJ+2glXk/4fWRCLVhHDvN60UnPl8mUBx
6OoYsipgs+FiyZr3ZKwFZcxwTzFdJX6jFYASaT66+KT8mAUYNMRrCa57U/BNK0NerPkKtWe3JUQt
glxXoYLW2Hw3yxprrDaAvLWBFfPl7UdyGybFnU9PNJ7Y+FJVYRti2qDnxXslIgh0aQQT7YhnOoX1
znQ1yEiFzzfbv7jq9cSYFlq6tufCr/PTa7XVNyEizovP7168cHCc74ouMZKSS9Q9ftuR77GzerHL
5s3vD+3/8vJIvpK+6yczXgpbnZe0TZShY2g2pTW41oeywAfoDh2OOI7+mP5AA3FMSHmrpPlo5orl
o3Yop2fHwieIH4b6cbmZETVXBLAXL7gjSY2oLV/Mx+pe+oPMaokDtDwjMT5dUHI2UrmReIuSESCt
/f34r8ZwNKnKbxcjAlOkv9gQP5HyauboDJ3G2XBvmRlhaztiSvyxrrIGm3XtxGIEhGDqU8TD1T9i
uabp5G2iQKnxRtbqVlOkuXxB8luyzRfwHOBLZS8CrK3t82eCsqpUQUcF17Bs5MwT9Qm11miCgyCB
GUAmHzhtIxk/l3CcQyL/QEIrgQkZ8ygT3RNbOqqYGvnoK1ZPVitM84R8SRpSNmpIB52ytNxCg3rG
ujPYHCvZWKJmaSCbnTVnurvJkQDYTUVM7uZ9KMQIt+G3zNIW/hzvYSCEWxjL4mfU4A28L17620xo
Oxc7/NBqu6tnUXfntleM78ikpA1xvH/c0DeQOzsvqiyeWKVphHkYLpVYsiVKOwdO4qPBDhn6sAFb
Cn0TOgy2vI9j4KIYdG7jCjPJBL6ywueAOydk8AiLiFis2aD9BXplzVnfcwRQQFFVWofV+NVtlPJv
U4R9ttukhwx+fubjWpFrs1ub+F0DW1K/ckjowpwLc/7PWd5fE6kdYPa5CKrmYB/1weCwMlL/ARio
6KqVaLBwyECznDFWPHBUk/MWEwW/EpxpDGe1zNH41ofaFcfjzm8+djPzAHK3kRkZ3+vnpQHoI2rb
jBmoW1P+nbhdIAIy+2WShZ5E/0TkdkesJ3SOwX0j6l1ZY2MrW8AeIke2pN606OsSopuTu/UPcNpq
fKyE+3lQsUy+/jLhCXSnrJWM9dOtMl7pEmjMzUV1rODnWbAJNPYNzRY8ZdsZ2CVEq6JHicjQcJuS
OK6m81Jy+AF0A0wEUpbtcMUgRKzJdWiiMPHZy5e/m9uQA/tCL6txPYiVx8YrxLA1FZWLszvAnDvP
/crp/tYMhfP+FtB02wqkNW3FeCja7xVWL+E+8TzDfEwpkl8yC4tIAD2YPe2GI0DveEnnIq/r5tr1
sXgJsDaj3gVva9GA/mUJENf9wcFil0irGG86Rv1T4ViFK8IqSVn5ZPwwwY6PHrtKPJVW4En6ny1v
MtYsuP0Imuu07Amfh5SU3tt1QN0v9cM4utx84tr5av3DvnFQt0jFs8zkVaQsJOPK8DXKFL0WFOAk
s2vDYeN8zkF54Eo5At9J+XRVhqki6cd7GE1u5ZwXlEpOsuy9m//UCtFUzY+bsYqiBZxrBeLQNJay
K23AXxSle5RaMWveWRFNw5/wXIDO0Ilfgkh+7rSdHwFZsOSpNW97uyDaRJYn7AoO3x0Hh37/S/mV
uJd+X1FinS3iuMhwAldO1ZCUJ+F1rS8m2CUhwlm7pREaxBsn5V7I56Nk5r5WhauP7JM60JcSh5/j
HlmovWZCrbSr5OPMo7c1t6xM+4uvU63O/RC9w0iLHbBFnOjFHcylA2xQ1WWAydyj/Qoh6Obe0L1h
DUg5DXWJSIgSHiK5mu3I6mTuhiU2nCS5cvSDlHzLWBK3eI+uWVQVgzrD8mmgLwfvPl5T4YwRC5XJ
YftFgXgVCpClGbzTskVNv/LYHIuiKNPdfe+G9yWXykAaBgvFipugZTHcuaEAF6PWVg2U8OjE9iQA
NVJKdaZ2gKGG77cR/Wvfq3plV3F+ysZo6tsMce6WSdGf1fuU2SZmFvAneXH6xemRFKnyIUx4+uD5
qrWbc0kmRDRMzm4PSqwJT010QM77QL8gCgGH/D2Pm944YIdU3LSr74Zs4+f+IV54moPEmAP58tmy
fmRNVLXbQ9WVvsJcJLAk7nnc0CETfB7on/mZ4nv1976V+scNg3VEBYMFwIH9tgulp2CrTsquT3Se
l4wO3sSdTG+V9TeA/2IyjRLgwOWCIqbHoXAoClkJaZy2Lc6wK4l55Wlp42Uxhs+nSjN5xK780pdE
XOZswda0WL+0snRYp93CmiL/MJKl9OSk3K2bCDE5xz7L7/zprAw2fj8G70BNpKloCbY3wZnZnSIE
dVfEXPOfhqVMw/OE9g8WGtifoQUrAP1Lw2LOEAVCoq3y8LsX+Agvetg/ocR2AF0Cel/nbznu3MFt
eNzaMsRxji67hk6a/lNY8ETEmiDb6UBK2ijGEoIjajPBEa+YQD/JqO/y+1onirNEqiluW1UTafFu
BefzQ/SaDPYCnDFfsOywyvhsxKIInkcOYKTgL5v8+PkYJxbIaSv1S7+fo4Fm5i4jGRbBOd8Xt0dM
H7OZZb4X8YfIR/wTkYm7K1b741hqfex4cB8VI4PQSZD07aU92zWMvNNS1mhpd8NzsPOHHUeakKbe
bkt4eClatjqsi3LDeYYV2XY7x9TlxUUqcD0+1zmM9lfa+hkjKZTNpmsZ6g0ZWACUBlwNKEo6Tqmy
rtiEHEqTigxC9Oo3PU7/Uv9fbWNJyL5RgWtWX4plL/HDwUYbNDKSPx3LuK7pWRbodyReOBTTKiBp
SaPwB7u3VUM1KygrORs4ssVy+L6bOwCeyWHD+R8jC577Aiylq1K4t0lXybqQ0A1TIY/qCYFCop5X
b0wXa9UvIEA2N5bYPPBogLJ70Tr8a9fJDHvr6RavJlRQnJF+76C7eonf26GeB3JgOkklkHmTjCf3
GlNaEEfI7oH4u0NtCuWNivAnbEMn+LEP2672IaGRPi0NNlskF6DOODxy8OvulFw6Npu5lpY2hN89
/KgyIRyXhVHvn26udHcIgBuU/jZb07FbOGdziuS8Gqe9DsmVT04sP0wUL1m3xKdoC2mRVxbOe7qP
i92PoSRzlpJBhsuymfMETDM7a9PkQajYEJ26SXasANqx9XZ/3eZCeK7OfD6gtecayfBrtCHMCHCK
HQv8Ak9ZCo3+ExD34GBJXd7S1hMRAv9cm1TdCahNvTXld7Rlq78b1liZ4rHfh3w880wAFdc/hbNJ
LRZas0AQbbbRIIG6XQc+dqUqzUm5Go2m3hXzab2VLaOQvBb9BklvqEX3JqIxCZovZc0vvWdJUQOf
l8l6Oy5JdbuYRri1kiYh6Qxhk+kwijmrgesBjiSKUGBbuMB6jjmEAv0380QiGYCAUPkGArmBqyRt
Rj3W2Ng5Ar04DXUQWNYXARVftStqaEAqQaTto//Sk3i0HIfWkVOf7r7VDGcpTWc5efHwXuDrNt+0
fpAObUQZfUJ6Foh3QpnVeinSeospQWj2xh4Eq6XChXlWcS3Y92GCKzJDbASzbmCtMQJhaXEnULl3
GrOzIL1jtdPZQx+sfIu4flE+8IRlHTDFWJlimYCW6w7EK2105PU25yCnzg==
`protect end_protected
